VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_8
  CLASS BLOCK ;
  FOREIGN tt_um_test_8 ;
  ORIGIN 0.030 0.000 ;
  SIZE 151.740 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 142.830 224.760 143.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 145.590 224.760 145.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 140.070 224.760 140.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 52.520 142.525 53.115 142.865 ;
        RECT 52.520 141.205 52.695 142.525 ;
        RECT 52.520 141.100 53.115 141.205 ;
        RECT 52.520 140.800 53.900 141.100 ;
        RECT 52.520 140.655 53.115 140.800 ;
      LAYER mcon ;
        RECT 53.630 140.830 53.870 141.070 ;
      LAYER met1 ;
        RECT 53.570 140.800 118.730 141.100 ;
      LAYER via ;
        RECT 118.400 140.800 118.700 141.100 ;
      LAYER met2 ;
        RECT 118.400 83.300 118.700 141.130 ;
        RECT 118.410 83.265 118.690 83.300 ;
      LAYER via2 ;
        RECT 118.410 83.310 118.690 83.590 ;
      LAYER met3 ;
        RECT 118.385 83.600 118.715 83.615 ;
        RECT 118.385 83.300 147.900 83.600 ;
        RECT 118.385 83.285 118.715 83.300 ;
        RECT 147.600 4.000 147.900 83.300 ;
        RECT 147.600 3.700 151.400 4.000 ;
        RECT 151.100 0.980 151.400 3.700 ;
        RECT 150.800 0.020 151.700 0.980 ;
      LAYER via3 ;
        RECT 150.800 0.050 151.700 0.950 ;
      LAYER met4 ;
        RECT 150.810 0.955 151.710 1.000 ;
        RECT 150.795 0.045 151.710 0.955 ;
        RECT 150.810 0.000 151.710 0.045 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 29.520 159.700 29.850 159.715 ;
        RECT 28.350 159.500 29.850 159.700 ;
        RECT 29.520 159.475 29.850 159.500 ;
      LAYER mcon ;
        RECT 28.365 159.515 28.535 159.685 ;
      LAYER met1 ;
        RECT 23.470 159.700 23.730 159.760 ;
        RECT 16.950 159.500 23.730 159.700 ;
        RECT 16.950 135.500 17.250 159.500 ;
        RECT 23.470 159.440 23.730 159.500 ;
        RECT 25.570 159.700 25.830 159.760 ;
        RECT 28.305 159.700 28.595 159.715 ;
        RECT 25.570 159.500 28.595 159.700 ;
        RECT 25.570 159.440 25.830 159.500 ;
        RECT 28.305 159.485 28.595 159.500 ;
        RECT 16.950 135.200 82.080 135.500 ;
      LAYER via ;
        RECT 23.470 159.470 23.730 159.730 ;
        RECT 25.570 159.470 25.830 159.730 ;
        RECT 81.750 135.200 82.050 135.500 ;
      LAYER met2 ;
        RECT 23.440 159.700 23.760 159.730 ;
        RECT 25.540 159.700 25.860 159.730 ;
        RECT 23.440 159.500 25.860 159.700 ;
        RECT 23.440 159.470 23.760 159.500 ;
        RECT 25.540 159.470 25.860 159.500 ;
        RECT 81.750 78.450 82.050 135.530 ;
        RECT 81.760 78.415 82.040 78.450 ;
      LAYER via2 ;
        RECT 81.760 78.460 82.040 78.740 ;
      LAYER met3 ;
        RECT 81.735 78.750 82.065 78.765 ;
        RECT 81.735 78.450 127.750 78.750 ;
        RECT 81.735 78.435 82.065 78.450 ;
        RECT 127.450 1.950 127.750 78.450 ;
        RECT 127.450 1.650 132.100 1.950 ;
        RECT 131.800 0.980 132.100 1.650 ;
        RECT 131.500 0.020 132.400 0.980 ;
      LAYER via3 ;
        RECT 131.500 0.050 132.400 0.950 ;
      LAYER met4 ;
        RECT 131.490 0.955 132.390 1.000 ;
        RECT 131.490 0.045 132.405 0.955 ;
        RECT 131.490 0.000 132.390 0.045 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 31.020 173.850 31.350 173.865 ;
        RECT 30.000 173.650 31.350 173.850 ;
        RECT 31.020 173.625 31.350 173.650 ;
      LAYER mcon ;
        RECT 30.015 173.665 30.185 173.835 ;
      LAYER met1 ;
        RECT 29.955 173.850 30.245 173.865 ;
        RECT 13.750 173.650 30.245 173.850 ;
        RECT 13.750 131.550 14.050 173.650 ;
        RECT 29.955 173.635 30.245 173.650 ;
        RECT 13.750 131.250 76.780 131.550 ;
      LAYER via ;
        RECT 76.450 131.250 76.750 131.550 ;
      LAYER met2 ;
        RECT 76.450 73.600 76.750 131.580 ;
        RECT 76.460 73.565 76.740 73.600 ;
      LAYER via2 ;
        RECT 76.460 73.610 76.740 73.890 ;
      LAYER met3 ;
        RECT 76.435 73.900 76.765 73.915 ;
        RECT 76.435 73.600 108.900 73.900 ;
        RECT 76.435 73.585 76.765 73.600 ;
        RECT 108.600 3.600 108.900 73.600 ;
        RECT 108.600 3.300 110.250 3.600 ;
        RECT 109.950 1.700 110.250 3.300 ;
        RECT 109.950 1.400 112.750 1.700 ;
        RECT 112.450 1.030 112.750 1.400 ;
        RECT 112.150 0.070 113.050 1.030 ;
      LAYER via3 ;
        RECT 112.150 0.100 113.050 1.000 ;
      LAYER met4 ;
        RECT 112.145 1.000 113.055 1.005 ;
        RECT 112.145 0.095 113.070 1.000 ;
        RECT 112.170 0.000 113.070 0.095 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 92.850 0.000 93.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 73.530 0.000 74.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 54.210 0.000 55.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 34.890 0.000 35.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 15.570 0.000 16.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 137.310 224.760 137.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 134.550 224.760 134.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 131.790 224.760 132.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 129.030 224.760 129.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 126.270 224.760 126.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 123.510 224.760 123.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 120.750 224.760 121.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 117.990 224.760 118.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 115.230 224.760 115.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 112.470 224.760 112.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 109.710 224.760 110.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 106.950 224.760 107.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 104.190 224.760 104.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 101.430 224.760 101.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 98.670 224.760 98.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 95.910 224.760 96.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 48.990 224.760 49.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 46.230 224.760 46.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 43.470 224.760 43.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 40.710 224.760 41.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 37.950 224.760 38.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 35.190 224.760 35.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 32.430 224.760 32.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 29.670 224.760 29.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 71.070 224.760 71.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 68.310 224.760 68.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 65.550 224.760 65.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 62.790 224.760 63.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 60.030 224.760 60.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 57.270 224.760 57.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 54.510 224.760 54.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 51.750 224.760 52.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 93.150 224.760 93.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 90.390 224.760 90.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 87.630 224.760 87.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 84.870 224.760 85.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 82.110 224.760 82.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 79.350 224.760 79.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 76.590 224.760 76.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 73.830 224.760 74.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 30.510 175.450 33.550 175.460 ;
        RECT 30.510 173.855 35.290 175.450 ;
        RECT 33.530 173.845 35.290 173.855 ;
        RECT 38.110 172.160 41.150 172.460 ;
        RECT 38.110 170.855 42.900 172.160 ;
        RECT 41.130 170.555 42.900 170.855 ;
        RECT 30.060 170.150 32.650 170.160 ;
        RECT 30.060 168.555 34.190 170.150 ;
        RECT 32.630 168.545 34.190 168.555 ;
        RECT 49.500 163.800 54.400 163.850 ;
        RECT 49.500 162.245 56.190 163.800 ;
        RECT 54.330 162.195 56.190 162.245 ;
        RECT 31.630 161.310 33.340 161.350 ;
        RECT 29.010 159.745 33.340 161.310 ;
        RECT 29.010 159.705 31.750 159.745 ;
        RECT 38.860 158.800 41.900 158.810 ;
        RECT 38.860 157.205 43.590 158.800 ;
        RECT 41.880 157.195 43.590 157.205 ;
        RECT 29.050 154.845 33.190 156.450 ;
        RECT 36.450 145.350 39.050 145.400 ;
        RECT 26.530 145.160 28.190 145.200 ;
        RECT 22.160 143.595 28.190 145.160 ;
        RECT 36.450 143.795 40.540 145.350 ;
        RECT 38.880 143.745 40.540 143.795 ;
        RECT 22.160 143.555 26.550 143.595 ;
        RECT 50.710 143.300 54.800 143.310 ;
        RECT 50.710 141.705 56.540 143.300 ;
        RECT 54.780 141.695 56.540 141.705 ;
      LAYER li1 ;
        RECT 30.700 175.185 32.080 175.355 ;
        RECT 31.040 174.045 31.250 175.185 ;
        RECT 34.640 175.175 35.100 175.345 ;
        RECT 34.725 174.010 35.015 175.175 ;
        RECT 38.300 172.185 39.680 172.355 ;
        RECT 39.255 171.045 39.585 172.185 ;
        RECT 42.250 171.885 42.710 172.055 ;
        RECT 42.335 170.720 42.625 171.885 ;
        RECT 30.250 169.885 31.630 170.055 ;
        RECT 30.590 168.745 30.800 169.885 ;
        RECT 33.540 169.875 34.000 170.045 ;
        RECT 33.625 168.710 33.915 169.875 ;
        RECT 49.690 163.575 52.910 163.745 ;
        RECT 50.745 162.725 50.915 163.575 ;
        RECT 51.585 163.065 51.755 163.575 ;
        RECT 55.540 163.525 56.000 163.695 ;
        RECT 55.625 162.360 55.915 163.525 ;
        RECT 29.200 161.035 30.580 161.205 ;
        RECT 32.690 161.075 33.150 161.245 ;
        RECT 29.540 159.895 29.750 161.035 ;
        RECT 32.775 159.910 33.065 161.075 ;
        RECT 39.050 158.535 40.430 158.705 ;
        RECT 40.005 157.395 40.335 158.535 ;
        RECT 42.940 158.525 43.400 158.695 ;
        RECT 43.025 157.360 43.315 158.525 ;
        RECT 29.240 156.175 30.620 156.345 ;
        RECT 32.540 156.175 33.000 156.345 ;
        RECT 29.580 155.035 29.790 156.175 ;
        RECT 32.625 155.010 32.915 156.175 ;
        RECT 36.640 145.125 38.020 145.295 ;
        RECT 22.350 144.885 24.650 145.055 ;
        RECT 27.540 144.925 28.000 145.095 ;
        RECT 22.865 144.485 23.800 144.885 ;
        RECT 27.625 143.760 27.915 144.925 ;
        RECT 36.980 143.985 37.190 145.125 ;
        RECT 39.890 145.075 40.350 145.245 ;
        RECT 39.975 143.910 40.265 145.075 ;
        RECT 50.900 143.035 53.200 143.205 ;
        RECT 51.415 142.635 52.350 143.035 ;
        RECT 55.890 143.025 56.350 143.195 ;
        RECT 55.975 141.860 56.265 143.025 ;
      LAYER mcon ;
        RECT 30.845 175.185 31.015 175.355 ;
        RECT 31.305 175.185 31.475 175.355 ;
        RECT 31.765 175.185 31.935 175.355 ;
        RECT 34.785 175.175 34.955 175.345 ;
        RECT 38.445 172.185 38.615 172.355 ;
        RECT 38.905 172.185 39.075 172.355 ;
        RECT 39.365 172.185 39.535 172.355 ;
        RECT 42.395 171.885 42.565 172.055 ;
        RECT 30.395 169.885 30.565 170.055 ;
        RECT 30.855 169.885 31.025 170.055 ;
        RECT 31.315 169.885 31.485 170.055 ;
        RECT 33.685 169.875 33.855 170.045 ;
        RECT 49.835 163.575 50.005 163.745 ;
        RECT 50.295 163.575 50.465 163.745 ;
        RECT 50.755 163.575 50.925 163.745 ;
        RECT 51.215 163.575 51.385 163.745 ;
        RECT 51.675 163.575 51.845 163.745 ;
        RECT 52.135 163.575 52.305 163.745 ;
        RECT 52.595 163.575 52.765 163.745 ;
        RECT 55.685 163.525 55.855 163.695 ;
        RECT 29.345 161.035 29.515 161.205 ;
        RECT 29.805 161.035 29.975 161.205 ;
        RECT 30.265 161.035 30.435 161.205 ;
        RECT 32.835 161.075 33.005 161.245 ;
        RECT 39.195 158.535 39.365 158.705 ;
        RECT 39.655 158.535 39.825 158.705 ;
        RECT 40.115 158.535 40.285 158.705 ;
        RECT 43.085 158.525 43.255 158.695 ;
        RECT 29.385 156.175 29.555 156.345 ;
        RECT 29.845 156.175 30.015 156.345 ;
        RECT 30.305 156.175 30.475 156.345 ;
        RECT 32.685 156.175 32.855 156.345 ;
        RECT 36.785 145.125 36.955 145.295 ;
        RECT 37.245 145.125 37.415 145.295 ;
        RECT 37.705 145.125 37.875 145.295 ;
        RECT 22.495 144.885 22.665 145.055 ;
        RECT 22.955 144.885 23.125 145.055 ;
        RECT 23.415 144.885 23.585 145.055 ;
        RECT 23.875 144.885 24.045 145.055 ;
        RECT 24.335 144.885 24.505 145.055 ;
        RECT 27.685 144.925 27.855 145.095 ;
        RECT 40.035 145.075 40.205 145.245 ;
        RECT 51.045 143.035 51.215 143.205 ;
        RECT 51.505 143.035 51.675 143.205 ;
        RECT 51.965 143.035 52.135 143.205 ;
        RECT 52.425 143.035 52.595 143.205 ;
        RECT 52.885 143.035 53.055 143.205 ;
        RECT 56.035 143.025 56.205 143.195 ;
      LAYER met1 ;
        RECT 31.460 176.395 31.750 176.430 ;
        RECT 31.460 176.070 31.765 176.395 ;
        RECT 31.475 175.510 31.765 176.070 ;
        RECT 30.700 175.030 32.080 175.510 ;
        RECT 34.700 175.500 35.000 176.880 ;
        RECT 34.640 175.020 35.100 175.500 ;
        RECT 42.350 173.300 42.650 173.330 ;
        RECT 42.345 172.970 42.650 173.300 ;
        RECT 38.300 172.400 39.680 172.510 ;
        RECT 40.100 172.400 40.400 172.430 ;
        RECT 38.300 172.100 40.400 172.400 ;
        RECT 42.345 172.210 42.645 172.970 ;
        RECT 38.300 172.030 39.680 172.100 ;
        RECT 40.100 172.070 40.400 172.100 ;
        RECT 42.250 171.730 42.710 172.210 ;
        RECT 28.205 170.655 30.855 170.945 ;
        RECT 23.910 170.195 24.200 170.230 ;
        RECT 28.205 170.195 28.495 170.655 ;
        RECT 30.565 170.210 30.855 170.655 ;
        RECT 23.905 169.905 28.495 170.195 ;
        RECT 23.910 169.870 24.200 169.905 ;
        RECT 30.250 169.730 31.630 170.210 ;
        RECT 33.600 170.200 33.895 170.880 ;
        RECT 33.540 169.720 34.000 170.200 ;
        RECT 54.750 164.895 55.900 164.900 ;
        RECT 51.385 164.605 55.900 164.895 ;
        RECT 51.385 163.900 51.675 164.605 ;
        RECT 53.620 164.600 53.980 164.605 ;
        RECT 54.750 164.595 55.900 164.605 ;
        RECT 49.690 163.420 52.910 163.900 ;
        RECT 55.595 163.850 55.900 164.595 ;
        RECT 55.540 163.370 56.000 163.850 ;
        RECT 29.510 162.345 29.800 162.380 ;
        RECT 29.510 162.020 29.805 162.345 ;
        RECT 33.600 162.145 33.895 162.180 ;
        RECT 29.515 161.360 29.805 162.020 ;
        RECT 32.750 161.850 33.895 162.145 ;
        RECT 32.750 161.400 33.045 161.850 ;
        RECT 33.600 161.820 33.895 161.850 ;
        RECT 29.200 160.880 30.580 161.360 ;
        RECT 32.690 160.920 33.150 161.400 ;
        RECT 43.000 159.900 43.300 159.930 ;
        RECT 39.500 159.895 43.300 159.900 ;
        RECT 39.365 159.600 43.300 159.895 ;
        RECT 39.365 158.860 39.655 159.600 ;
        RECT 39.050 158.380 40.430 158.860 ;
        RECT 43.000 158.850 43.300 159.600 ;
        RECT 42.940 158.370 43.400 158.850 ;
        RECT 33.500 156.800 33.800 156.830 ;
        RECT 28.060 156.500 28.350 156.530 ;
        RECT 32.650 156.500 33.800 156.800 ;
        RECT 28.055 156.210 30.620 156.500 ;
        RECT 28.060 156.170 28.350 156.210 ;
        RECT 29.240 156.020 30.620 156.210 ;
        RECT 32.540 156.020 33.000 156.500 ;
        RECT 33.500 156.470 33.800 156.500 ;
        RECT 37.720 146.400 38.085 146.405 ;
        RECT 37.000 146.395 40.250 146.400 ;
        RECT 36.955 146.095 40.250 146.395 ;
        RECT 27.650 146.000 27.955 146.035 ;
        RECT 27.645 145.995 27.955 146.000 ;
        RECT 23.125 145.705 27.955 145.995 ;
        RECT 23.125 145.210 23.415 145.705 ;
        RECT 27.645 145.670 27.955 145.705 ;
        RECT 27.645 145.250 27.950 145.670 ;
        RECT 36.955 145.450 37.245 146.095 ;
        RECT 22.350 144.730 24.650 145.210 ;
        RECT 27.540 144.770 28.000 145.250 ;
        RECT 36.640 144.970 38.020 145.450 ;
        RECT 39.945 145.400 40.250 146.095 ;
        RECT 39.890 144.920 40.350 145.400 ;
        RECT 52.150 144.345 52.440 144.380 ;
        RECT 52.135 144.020 52.440 144.345 ;
        RECT 52.135 143.360 52.425 144.020 ;
        RECT 50.900 142.880 53.200 143.360 ;
        RECT 55.950 143.350 56.250 144.380 ;
        RECT 55.890 142.870 56.350 143.350 ;
      LAYER via ;
        RECT 34.700 176.550 35.000 176.850 ;
        RECT 31.460 176.100 31.750 176.400 ;
        RECT 42.350 173.000 42.650 173.300 ;
        RECT 40.100 172.100 40.400 172.400 ;
        RECT 23.910 169.900 24.200 170.200 ;
        RECT 33.600 170.550 33.895 170.850 ;
        RECT 53.650 164.600 53.950 164.890 ;
        RECT 29.510 162.050 29.800 162.350 ;
        RECT 33.600 161.850 33.895 162.150 ;
        RECT 43.000 159.600 43.300 159.900 ;
        RECT 33.500 156.500 33.800 156.800 ;
        RECT 28.060 156.200 28.350 156.500 ;
        RECT 37.750 146.100 38.055 146.405 ;
        RECT 27.650 145.700 27.955 146.005 ;
        RECT 52.150 144.050 52.440 144.350 ;
        RECT 55.950 144.050 56.250 144.350 ;
      LAYER met2 ;
        RECT 34.060 176.850 34.340 176.885 ;
        RECT 34.050 176.550 35.030 176.850 ;
        RECT 34.060 176.515 34.340 176.550 ;
        RECT 30.760 176.400 31.040 176.435 ;
        RECT 30.750 176.100 31.780 176.400 ;
        RECT 30.760 176.065 31.040 176.100 ;
        RECT 41.510 173.300 41.790 173.335 ;
        RECT 41.500 173.000 42.680 173.300 ;
        RECT 41.510 172.965 41.790 173.000 ;
        RECT 41.010 172.400 41.290 172.435 ;
        RECT 40.070 172.100 41.290 172.400 ;
        RECT 41.010 172.065 41.290 172.100 ;
        RECT 34.560 170.850 34.840 170.885 ;
        RECT 33.570 170.550 34.850 170.850 ;
        RECT 34.560 170.515 34.840 170.550 ;
        RECT 17.960 170.200 18.240 170.235 ;
        RECT 17.950 169.900 24.230 170.200 ;
        RECT 17.960 169.865 18.240 169.900 ;
        RECT 53.650 165.790 53.950 165.800 ;
        RECT 53.615 165.510 53.985 165.790 ;
        RECT 53.650 164.570 53.950 165.510 ;
        RECT 28.760 162.350 29.040 162.385 ;
        RECT 28.750 162.050 29.830 162.350 ;
        RECT 33.570 162.140 34.950 162.150 ;
        RECT 28.760 162.015 29.040 162.050 ;
        RECT 33.570 161.860 34.985 162.140 ;
        RECT 33.570 161.850 34.950 161.860 ;
        RECT 42.970 159.890 44.200 159.900 ;
        RECT 42.970 159.610 44.235 159.890 ;
        RECT 42.970 159.600 44.200 159.610 ;
        RECT 33.470 156.790 34.650 156.800 ;
        RECT 33.470 156.510 34.685 156.790 ;
        RECT 33.470 156.500 34.650 156.510 ;
        RECT 26.900 156.490 28.380 156.500 ;
        RECT 26.865 156.210 28.380 156.490 ;
        RECT 26.900 156.200 28.380 156.210 ;
        RECT 37.760 147.400 38.040 147.435 ;
        RECT 37.750 146.435 38.050 147.400 ;
        RECT 37.750 146.070 38.055 146.435 ;
        RECT 27.620 146.000 27.985 146.005 ;
        RECT 27.620 145.990 29.000 146.000 ;
        RECT 27.620 145.710 29.035 145.990 ;
        RECT 27.620 145.700 29.000 145.710 ;
        RECT 52.120 144.050 56.280 144.350 ;
      LAYER via2 ;
        RECT 34.060 176.560 34.340 176.840 ;
        RECT 30.760 176.110 31.040 176.390 ;
        RECT 41.510 173.010 41.790 173.290 ;
        RECT 41.010 172.110 41.290 172.390 ;
        RECT 34.560 170.560 34.840 170.840 ;
        RECT 17.960 169.910 18.240 170.190 ;
        RECT 20.060 169.910 20.340 170.190 ;
        RECT 53.660 165.510 53.940 165.790 ;
        RECT 28.760 162.060 29.040 162.340 ;
        RECT 34.660 161.860 34.940 162.140 ;
        RECT 43.910 159.610 44.190 159.890 ;
        RECT 34.360 156.510 34.640 156.790 ;
        RECT 26.910 156.210 27.190 156.490 ;
        RECT 37.760 147.110 38.040 147.390 ;
        RECT 28.710 145.710 28.990 145.990 ;
        RECT 54.860 144.060 55.140 144.340 ;
      LAYER met3 ;
        RECT 30.650 179.100 36.750 179.400 ;
        RECT 30.650 177.750 30.950 179.100 ;
        RECT 29.250 177.450 32.850 177.750 ;
        RECT 29.250 176.400 29.550 177.450 ;
        RECT 32.550 176.850 32.850 177.450 ;
        RECT 34.035 176.850 34.365 176.865 ;
        RECT 32.550 176.550 34.365 176.850 ;
        RECT 34.035 176.535 34.365 176.550 ;
        RECT 30.735 176.400 31.065 176.415 ;
        RECT 20.050 176.100 31.065 176.400 ;
        RECT -0.030 170.200 2.030 171.050 ;
        RECT 5.810 170.200 6.190 170.210 ;
        RECT -0.030 169.900 6.190 170.200 ;
        RECT -0.030 169.050 2.030 169.900 ;
        RECT 5.810 169.890 6.190 169.900 ;
        RECT 11.090 170.200 11.410 170.240 ;
        RECT 20.050 170.215 20.350 176.100 ;
        RECT 30.735 176.085 31.065 176.100 ;
        RECT 36.450 175.050 36.750 179.100 ;
        RECT 36.450 174.750 40.950 175.050 ;
        RECT 36.450 172.200 36.750 174.750 ;
        RECT 40.650 174.500 40.950 174.750 ;
        RECT 40.650 174.200 43.600 174.500 ;
        RECT 40.650 173.300 40.950 174.200 ;
        RECT 41.485 173.300 41.815 173.315 ;
        RECT 40.650 173.000 41.815 173.300 ;
        RECT 41.485 172.985 41.815 173.000 ;
        RECT 35.200 171.900 36.750 172.200 ;
        RECT 40.985 172.400 41.315 172.415 ;
        RECT 43.300 172.400 43.600 174.200 ;
        RECT 40.985 172.100 43.600 172.400 ;
        RECT 40.985 172.085 41.315 172.100 ;
        RECT 34.535 170.850 34.865 170.865 ;
        RECT 35.200 170.850 35.500 171.900 ;
        RECT 34.535 170.550 35.500 170.850 ;
        RECT 34.535 170.535 34.865 170.550 ;
        RECT 17.935 170.200 18.265 170.215 ;
        RECT 11.090 169.900 18.265 170.200 ;
        RECT 11.090 169.860 11.410 169.900 ;
        RECT 15.750 168.500 16.050 169.900 ;
        RECT 17.935 169.885 18.265 169.900 ;
        RECT 20.035 169.885 20.365 170.215 ;
        RECT 15.750 168.200 23.200 168.500 ;
        RECT 22.900 162.350 23.200 168.200 ;
        RECT 41.750 166.850 53.950 167.150 ;
        RECT 41.750 163.200 42.050 166.850 ;
        RECT 53.650 165.815 53.950 166.850 ;
        RECT 53.635 165.485 53.965 165.815 ;
        RECT 27.950 162.900 44.200 163.200 ;
        RECT 27.950 162.350 28.250 162.900 ;
        RECT 28.735 162.350 29.065 162.365 ;
        RECT 22.900 162.050 29.065 162.350 ;
        RECT 34.650 162.165 34.950 162.900 ;
        RECT 26.900 157.400 27.200 162.050 ;
        RECT 28.735 162.035 29.065 162.050 ;
        RECT 34.635 161.835 34.965 162.165 ;
        RECT 43.900 159.915 44.200 162.900 ;
        RECT 43.885 159.585 44.215 159.915 ;
        RECT 29.900 157.550 34.650 157.850 ;
        RECT 29.900 157.400 30.200 157.550 ;
        RECT 25.550 157.100 30.200 157.400 ;
        RECT 25.550 149.150 25.850 157.100 ;
        RECT 26.900 156.515 27.200 157.100 ;
        RECT 34.350 156.815 34.650 157.550 ;
        RECT 26.885 156.185 27.215 156.515 ;
        RECT 34.335 156.485 34.665 156.815 ;
        RECT 30.950 151.100 43.450 151.400 ;
        RECT 30.950 149.150 31.250 151.100 ;
        RECT 25.550 148.850 32.800 149.150 ;
        RECT 25.550 147.200 25.850 148.850 ;
        RECT 32.500 147.400 32.800 148.850 ;
        RECT 37.735 147.400 38.065 147.415 ;
        RECT 25.550 146.900 29.000 147.200 ;
        RECT 32.500 147.100 38.065 147.400 ;
        RECT 37.735 147.085 38.065 147.100 ;
        RECT 28.700 146.015 29.000 146.900 ;
        RECT 43.150 146.750 43.450 151.100 ;
        RECT 43.150 146.450 55.150 146.750 ;
        RECT 28.685 145.685 29.015 146.015 ;
        RECT 54.850 144.365 55.150 146.450 ;
        RECT 54.835 144.035 55.165 144.365 ;
      LAYER via3 ;
        RECT 0.000 169.050 2.000 171.050 ;
        RECT 5.840 169.890 6.160 170.210 ;
        RECT 11.090 169.890 11.410 170.210 ;
      LAYER met4 ;
        RECT 0.000 171.055 2.000 220.760 ;
        RECT -0.005 169.045 2.005 171.055 ;
        RECT 5.835 170.200 6.165 170.215 ;
        RECT 11.085 170.200 11.415 170.215 ;
        RECT 5.835 169.900 11.415 170.200 ;
        RECT 5.835 169.885 6.165 169.900 ;
        RECT 11.085 169.885 11.415 169.900 ;
        RECT 0.000 5.000 2.000 169.045 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 34.785 172.860 34.955 173.385 ;
        RECT 42.395 169.570 42.565 170.095 ;
        RECT 33.685 167.560 33.855 168.085 ;
        RECT 55.685 161.210 55.855 161.735 ;
        RECT 32.835 158.760 33.005 159.285 ;
        RECT 43.085 156.210 43.255 156.735 ;
        RECT 32.685 153.860 32.855 154.385 ;
        RECT 27.685 142.610 27.855 143.135 ;
        RECT 40.035 142.760 40.205 143.285 ;
        RECT 56.035 140.710 56.205 141.235 ;
      LAYER li1 ;
        RECT 31.020 172.635 31.250 173.455 ;
        RECT 30.700 172.465 32.080 172.635 ;
        RECT 34.725 172.625 35.015 173.350 ;
        RECT 34.640 172.455 35.100 172.625 ;
        RECT 38.405 169.635 38.645 170.445 ;
        RECT 39.315 169.635 39.585 170.445 ;
        RECT 38.300 169.465 39.680 169.635 ;
        RECT 42.335 169.335 42.625 170.060 ;
        RECT 42.250 169.165 42.710 169.335 ;
        RECT 30.570 167.335 30.800 168.155 ;
        RECT 30.250 167.165 31.630 167.335 ;
        RECT 33.625 167.325 33.915 168.050 ;
        RECT 33.540 167.155 34.000 167.325 ;
        RECT 49.825 161.025 50.155 161.415 ;
        RECT 50.665 161.025 50.995 161.415 ;
        RECT 52.535 161.025 52.825 161.860 ;
        RECT 49.690 160.855 52.910 161.025 ;
        RECT 55.625 160.975 55.915 161.700 ;
        RECT 55.540 160.805 56.000 160.975 ;
        RECT 29.520 158.485 29.750 159.305 ;
        RECT 32.775 158.525 33.065 159.250 ;
        RECT 29.200 158.315 30.580 158.485 ;
        RECT 32.690 158.355 33.150 158.525 ;
        RECT 39.155 155.985 39.395 156.795 ;
        RECT 40.065 155.985 40.335 156.795 ;
        RECT 39.050 155.815 40.430 155.985 ;
        RECT 43.025 155.975 43.315 156.700 ;
        RECT 42.940 155.805 43.400 155.975 ;
        RECT 29.560 153.625 29.790 154.445 ;
        RECT 32.625 153.625 32.915 154.350 ;
        RECT 29.240 153.455 30.620 153.625 ;
        RECT 32.540 153.455 33.000 153.625 ;
        RECT 22.865 142.335 23.800 142.735 ;
        RECT 27.625 142.375 27.915 143.100 ;
        RECT 36.960 142.575 37.190 143.395 ;
        RECT 36.640 142.405 38.020 142.575 ;
        RECT 39.975 142.525 40.265 143.250 ;
        RECT 22.350 142.165 24.650 142.335 ;
        RECT 27.540 142.205 28.000 142.375 ;
        RECT 39.890 142.355 40.350 142.525 ;
        RECT 51.415 140.485 52.350 140.885 ;
        RECT 50.900 140.315 53.200 140.485 ;
        RECT 55.975 140.475 56.265 141.200 ;
        RECT 55.890 140.305 56.350 140.475 ;
      LAYER mcon ;
        RECT 30.845 172.465 31.015 172.635 ;
        RECT 31.305 172.465 31.475 172.635 ;
        RECT 31.765 172.465 31.935 172.635 ;
        RECT 34.785 172.455 34.955 172.625 ;
        RECT 38.445 169.465 38.615 169.635 ;
        RECT 38.905 169.465 39.075 169.635 ;
        RECT 39.365 169.465 39.535 169.635 ;
        RECT 42.395 169.165 42.565 169.335 ;
        RECT 30.395 167.165 30.565 167.335 ;
        RECT 30.855 167.165 31.025 167.335 ;
        RECT 31.315 167.165 31.485 167.335 ;
        RECT 33.685 167.155 33.855 167.325 ;
        RECT 49.835 160.855 50.005 161.025 ;
        RECT 50.295 160.855 50.465 161.025 ;
        RECT 50.755 160.855 50.925 161.025 ;
        RECT 51.215 160.855 51.385 161.025 ;
        RECT 51.675 160.855 51.845 161.025 ;
        RECT 52.135 160.855 52.305 161.025 ;
        RECT 52.595 160.855 52.765 161.025 ;
        RECT 55.685 160.805 55.855 160.975 ;
        RECT 29.345 158.315 29.515 158.485 ;
        RECT 29.805 158.315 29.975 158.485 ;
        RECT 30.265 158.315 30.435 158.485 ;
        RECT 32.835 158.355 33.005 158.525 ;
        RECT 39.195 155.815 39.365 155.985 ;
        RECT 39.655 155.815 39.825 155.985 ;
        RECT 40.115 155.815 40.285 155.985 ;
        RECT 43.085 155.805 43.255 155.975 ;
        RECT 29.385 153.455 29.555 153.625 ;
        RECT 29.845 153.455 30.015 153.625 ;
        RECT 30.305 153.455 30.475 153.625 ;
        RECT 32.685 153.455 32.855 153.625 ;
        RECT 36.785 142.405 36.955 142.575 ;
        RECT 37.245 142.405 37.415 142.575 ;
        RECT 37.705 142.405 37.875 142.575 ;
        RECT 22.495 142.165 22.665 142.335 ;
        RECT 22.955 142.165 23.125 142.335 ;
        RECT 23.415 142.165 23.585 142.335 ;
        RECT 23.875 142.165 24.045 142.335 ;
        RECT 24.335 142.165 24.505 142.335 ;
        RECT 27.685 142.205 27.855 142.375 ;
        RECT 40.035 142.355 40.205 142.525 ;
        RECT 51.045 140.315 51.215 140.485 ;
        RECT 51.505 140.315 51.675 140.485 ;
        RECT 51.965 140.315 52.135 140.485 ;
        RECT 52.425 140.315 52.595 140.485 ;
        RECT 52.885 140.315 53.055 140.485 ;
        RECT 56.035 140.305 56.205 140.475 ;
      LAYER met1 ;
        RECT 30.700 172.310 32.080 172.790 ;
        RECT 23.860 172.045 24.150 172.080 ;
        RECT 31.015 172.045 31.305 172.310 ;
        RECT 34.640 172.300 35.100 172.780 ;
        RECT 23.855 171.755 31.305 172.045 ;
        RECT 34.750 171.770 35.050 172.300 ;
        RECT 23.860 171.720 24.150 171.755 ;
        RECT 37.660 169.600 37.950 169.630 ;
        RECT 38.300 169.600 39.680 169.790 ;
        RECT 37.655 169.310 39.680 169.600 ;
        RECT 37.660 169.270 37.950 169.310 ;
        RECT 42.250 169.010 42.710 169.490 ;
        RECT 42.300 168.270 42.600 169.010 ;
        RECT 30.250 167.010 31.630 167.490 ;
        RECT 25.660 166.495 25.950 166.530 ;
        RECT 30.565 166.495 30.855 167.010 ;
        RECT 33.540 167.000 34.000 167.480 ;
        RECT 25.655 166.205 30.855 166.495 ;
        RECT 33.595 166.680 33.895 167.000 ;
        RECT 33.595 166.350 33.900 166.680 ;
        RECT 33.600 166.320 33.900 166.350 ;
        RECT 25.660 166.170 25.950 166.205 ;
        RECT 48.760 160.990 49.050 161.030 ;
        RECT 49.690 160.990 52.910 161.180 ;
        RECT 48.755 160.700 52.910 160.990 ;
        RECT 48.760 160.670 49.050 160.700 ;
        RECT 55.540 160.650 56.000 161.130 ;
        RECT 55.600 159.720 55.900 160.650 ;
        RECT 29.200 158.160 30.580 158.640 ;
        RECT 32.690 158.250 33.150 158.680 ;
        RECT 33.600 158.250 33.900 158.280 ;
        RECT 32.690 158.200 33.900 158.250 ;
        RECT 25.560 157.845 25.850 157.880 ;
        RECT 29.515 157.845 29.805 158.160 ;
        RECT 32.745 157.950 33.900 158.200 ;
        RECT 33.600 157.920 33.900 157.950 ;
        RECT 25.555 157.555 29.805 157.845 ;
        RECT 25.560 157.520 25.850 157.555 ;
        RECT 38.260 155.950 38.550 155.980 ;
        RECT 39.050 155.950 40.430 156.140 ;
        RECT 38.255 155.660 40.430 155.950 ;
        RECT 38.260 155.620 38.550 155.660 ;
        RECT 42.940 155.650 43.400 156.130 ;
        RECT 43.045 155.085 43.350 155.650 ;
        RECT 43.045 154.750 43.355 155.085 ;
        RECT 43.050 154.720 43.355 154.750 ;
        RECT 29.240 153.300 30.620 153.780 ;
        RECT 32.540 153.300 33.000 153.780 ;
        RECT 29.555 153.130 29.845 153.300 ;
        RECT 29.555 152.805 29.850 153.130 ;
        RECT 29.560 152.770 29.850 152.805 ;
        RECT 32.600 152.600 32.900 153.300 ;
        RECT 32.570 152.300 32.930 152.600 ;
        RECT 35.860 142.540 36.150 142.580 ;
        RECT 36.640 142.540 38.020 142.730 ;
        RECT 22.350 142.010 24.650 142.490 ;
        RECT 27.540 142.050 28.000 142.530 ;
        RECT 35.855 142.250 38.020 142.540 ;
        RECT 35.860 142.220 36.150 142.250 ;
        RECT 39.890 142.200 40.350 142.680 ;
        RECT 28.450 142.050 28.750 142.080 ;
        RECT 23.125 141.780 23.415 142.010 ;
        RECT 23.110 141.455 23.415 141.780 ;
        RECT 27.600 141.750 28.750 142.050 ;
        RECT 39.950 141.950 40.250 142.200 ;
        RECT 28.450 141.720 28.750 141.750 ;
        RECT 39.955 141.700 40.250 141.950 ;
        RECT 23.110 141.420 23.400 141.455 ;
        RECT 39.920 141.405 40.280 141.700 ;
        RECT 50.210 140.450 50.500 140.480 ;
        RECT 50.900 140.450 53.200 140.640 ;
        RECT 50.205 140.160 53.200 140.450 ;
        RECT 50.210 140.120 50.500 140.160 ;
        RECT 55.890 140.150 56.350 140.630 ;
        RECT 55.950 139.420 56.250 140.150 ;
      LAYER via ;
        RECT 23.860 171.750 24.150 172.050 ;
        RECT 34.750 171.800 35.050 172.100 ;
        RECT 37.660 169.300 37.950 169.600 ;
        RECT 42.300 168.300 42.600 168.600 ;
        RECT 25.660 166.200 25.950 166.500 ;
        RECT 33.600 166.350 33.900 166.650 ;
        RECT 48.760 160.700 49.050 161.000 ;
        RECT 55.600 159.750 55.900 160.050 ;
        RECT 25.560 157.550 25.850 157.850 ;
        RECT 33.600 157.950 33.900 158.250 ;
        RECT 38.260 155.650 38.550 155.950 ;
        RECT 43.050 154.750 43.355 155.055 ;
        RECT 29.560 152.800 29.850 153.100 ;
        RECT 32.600 152.300 32.900 152.600 ;
        RECT 35.860 142.250 36.150 142.550 ;
        RECT 28.450 141.750 28.750 142.050 ;
        RECT 23.110 141.450 23.400 141.750 ;
        RECT 39.950 141.405 40.250 141.700 ;
        RECT 50.210 140.150 50.500 140.450 ;
        RECT 55.950 139.450 56.250 139.750 ;
      LAYER met2 ;
        RECT 17.960 172.050 18.240 172.085 ;
        RECT 17.950 171.750 24.180 172.050 ;
        RECT 31.550 171.800 35.080 172.100 ;
        RECT 17.960 171.715 18.240 171.750 ;
        RECT 31.550 166.650 31.850 171.800 ;
        RECT 35.700 169.300 37.980 169.600 ;
        RECT 35.700 168.600 36.000 169.300 ;
        RECT 35.700 168.300 42.630 168.600 ;
        RECT 19.060 166.500 19.340 166.535 ;
        RECT 19.050 166.200 25.980 166.500 ;
        RECT 31.550 166.350 33.930 166.650 ;
        RECT 19.060 166.165 19.340 166.200 ;
        RECT 21.000 164.300 21.300 166.200 ;
        RECT 31.550 164.300 31.850 166.350 ;
        RECT 35.700 164.300 36.000 168.300 ;
        RECT 21.000 164.000 36.000 164.300 ;
        RECT 21.000 157.850 21.300 164.000 ;
        RECT 35.700 161.000 36.000 164.000 ;
        RECT 35.700 160.700 49.080 161.000 ;
        RECT 35.700 158.250 36.000 160.700 ;
        RECT 47.200 160.050 47.500 160.700 ;
        RECT 47.200 159.750 55.930 160.050 ;
        RECT 33.570 157.950 36.000 158.250 ;
        RECT 21.000 157.550 25.880 157.850 ;
        RECT 21.000 153.100 21.300 157.550 ;
        RECT 35.700 155.950 36.000 157.950 ;
        RECT 35.700 155.650 38.580 155.950 ;
        RECT 37.400 155.050 37.700 155.650 ;
        RECT 43.020 155.050 43.385 155.055 ;
        RECT 37.400 154.750 43.385 155.050 ;
        RECT 21.000 152.800 29.880 153.100 ;
        RECT 21.000 141.750 21.300 152.800 ;
        RECT 28.700 151.750 29.000 152.800 ;
        RECT 32.600 151.750 32.900 152.630 ;
        RECT 28.700 151.450 32.900 151.750 ;
        RECT 31.100 142.250 36.180 142.550 ;
        RECT 31.100 142.050 31.400 142.250 ;
        RECT 28.420 141.750 31.400 142.050 ;
        RECT 21.000 141.450 23.430 141.750 ;
        RECT 21.000 139.500 21.300 141.450 ;
        RECT 31.100 140.450 31.400 141.750 ;
        RECT 39.950 140.450 40.250 141.730 ;
        RECT 31.100 140.150 50.530 140.450 ;
        RECT 31.100 139.500 31.400 140.150 ;
        RECT 21.000 139.200 31.400 139.500 ;
        RECT 49.500 138.950 49.800 140.150 ;
        RECT 54.800 139.450 56.280 139.750 ;
        RECT 54.800 138.950 55.100 139.450 ;
        RECT 49.500 138.650 55.100 138.950 ;
      LAYER via2 ;
        RECT 17.960 171.760 18.240 172.040 ;
        RECT 19.060 166.210 19.340 166.490 ;
      LAYER met3 ;
        RECT 17.935 172.050 18.265 172.065 ;
        RECT 9.550 171.750 18.265 172.050 ;
        RECT 9.550 168.150 9.850 171.750 ;
        RECT 17.935 171.735 18.265 171.750 ;
        RECT 9.550 167.850 13.050 168.150 ;
        RECT 2.970 166.500 5.030 167.350 ;
        RECT 12.750 166.500 13.050 167.850 ;
        RECT 19.035 166.500 19.365 166.515 ;
        RECT 2.970 166.200 19.365 166.500 ;
        RECT 2.970 165.350 5.030 166.200 ;
        RECT 19.035 166.185 19.365 166.200 ;
      LAYER via3 ;
        RECT 3.000 165.350 5.000 167.350 ;
      LAYER met4 ;
        RECT 3.000 167.355 5.000 220.760 ;
        RECT 2.995 165.345 5.005 167.355 ;
        RECT 3.000 5.000 5.000 165.345 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 30.845 172.465 31.015 172.635 ;
        RECT 38.450 169.465 38.620 169.635 ;
        RECT 30.395 167.165 30.565 167.335 ;
        RECT 49.835 160.855 50.005 161.025 ;
        RECT 29.345 158.315 29.515 158.485 ;
        RECT 39.200 155.815 39.370 155.985 ;
        RECT 29.385 153.455 29.555 153.625 ;
        RECT 36.785 142.405 36.955 142.575 ;
        RECT 22.500 142.165 22.670 142.335 ;
        RECT 51.050 140.315 51.220 140.485 ;
      LAYER li1 ;
        RECT 31.420 174.035 31.750 175.015 ;
        RECT 31.520 173.715 31.750 174.035 ;
        RECT 31.520 173.485 33.115 173.715 ;
        RECT 31.520 173.435 31.750 173.485 ;
        RECT 31.420 172.805 31.750 173.435 ;
        RECT 37.650 172.900 38.300 173.100 ;
        RECT 37.650 171.750 37.850 172.900 ;
        RECT 38.395 171.750 38.725 172.000 ;
        RECT 37.650 171.550 38.725 171.750 ;
        RECT 38.395 171.215 38.725 171.550 ;
        RECT 38.395 171.045 39.075 171.215 ;
        RECT 38.385 170.625 38.735 170.875 ;
        RECT 38.905 170.445 39.075 171.045 ;
        RECT 39.245 170.845 39.595 170.875 ;
        RECT 39.245 170.655 40.795 170.845 ;
        RECT 39.245 170.625 39.595 170.655 ;
        RECT 38.815 169.805 39.145 170.445 ;
        RECT 30.970 168.735 31.300 169.715 ;
        RECT 30.570 168.550 30.900 168.565 ;
        RECT 29.450 168.350 30.900 168.550 ;
        RECT 30.570 168.325 30.900 168.350 ;
        RECT 31.070 168.415 31.300 168.735 ;
        RECT 31.070 168.185 32.565 168.415 ;
        RECT 31.070 168.135 31.300 168.185 ;
        RECT 30.970 167.505 31.300 168.135 ;
        RECT 49.775 162.725 50.155 163.405 ;
        RECT 51.085 162.895 51.415 163.405 ;
        RECT 51.925 162.895 52.325 163.405 ;
        RECT 51.085 162.725 52.325 162.895 ;
        RECT 52.505 162.750 52.825 163.405 ;
        RECT 49.775 161.765 49.945 162.725 ;
        RECT 50.115 162.385 51.420 162.555 ;
        RECT 52.505 162.475 52.900 162.750 ;
        RECT 50.115 161.935 50.360 162.385 ;
        RECT 50.530 162.015 51.080 162.215 ;
        RECT 51.250 162.185 51.420 162.385 ;
        RECT 52.195 162.450 52.900 162.475 ;
        RECT 52.195 162.305 52.825 162.450 ;
        RECT 51.250 162.015 51.625 162.185 ;
        RECT 51.795 161.765 52.025 162.265 ;
        RECT 49.775 161.595 52.025 161.765 ;
        RECT 50.325 161.275 50.495 161.595 ;
        RECT 52.195 161.425 52.365 162.305 ;
        RECT 51.410 161.255 52.365 161.425 ;
        RECT 29.920 159.885 30.250 160.865 ;
        RECT 30.020 159.515 30.250 159.885 ;
        RECT 30.020 159.285 31.565 159.515 ;
        RECT 29.920 158.655 30.250 159.285 ;
        RECT 31.335 159.135 31.565 159.285 ;
        RECT 39.145 158.100 39.475 158.350 ;
        RECT 39.000 157.800 39.475 158.100 ;
        RECT 39.145 157.565 39.475 157.800 ;
        RECT 39.145 157.395 39.825 157.565 ;
        RECT 38.075 156.975 39.485 157.225 ;
        RECT 39.655 156.795 39.825 157.395 ;
        RECT 39.995 157.200 40.345 157.225 ;
        RECT 39.995 157.000 41.300 157.200 ;
        RECT 39.995 156.975 40.345 157.000 ;
        RECT 39.565 156.155 39.895 156.795 ;
        RECT 29.960 155.025 30.290 156.005 ;
        RECT 29.560 154.850 29.890 154.855 ;
        RECT 28.400 154.650 29.890 154.850 ;
        RECT 29.560 154.615 29.890 154.650 ;
        RECT 30.060 154.665 30.290 155.025 ;
        RECT 31.335 154.665 31.565 154.915 ;
        RECT 30.060 154.435 31.565 154.665 ;
        RECT 30.060 154.425 30.290 154.435 ;
        RECT 29.960 153.795 30.290 154.425 ;
        RECT 22.435 144.315 22.695 144.715 ;
        RECT 23.970 144.375 24.565 144.715 ;
        RECT 22.435 144.145 23.800 144.315 ;
        RECT 22.435 143.500 22.895 143.975 ;
        RECT 21.600 143.300 22.895 143.500 ;
        RECT 22.435 143.245 22.895 143.300 ;
        RECT 23.065 143.075 23.800 144.145 ;
        RECT 22.435 142.905 23.800 143.075 ;
        RECT 23.970 143.055 24.145 144.375 ;
        RECT 24.325 143.450 24.565 144.205 ;
        RECT 37.360 143.975 37.690 144.955 ;
        RECT 36.960 143.800 37.290 143.805 ;
        RECT 35.850 143.600 37.290 143.800 ;
        RECT 36.960 143.565 37.290 143.600 ;
        RECT 24.325 143.250 25.500 143.450 ;
        RECT 37.460 143.375 37.690 143.975 ;
        RECT 24.325 143.225 24.565 143.250 ;
        RECT 22.435 142.505 22.695 142.905 ;
        RECT 23.970 142.505 24.565 143.055 ;
        RECT 37.360 142.745 37.690 143.375 ;
        RECT 50.985 142.465 51.245 142.865 ;
        RECT 50.985 142.295 52.350 142.465 ;
        RECT 50.985 141.650 51.445 142.125 ;
        RECT 50.100 141.450 51.445 141.650 ;
        RECT 50.985 141.395 51.445 141.450 ;
        RECT 51.615 141.225 52.350 142.295 ;
        RECT 52.875 141.650 53.115 142.355 ;
        RECT 52.875 141.450 54.200 141.650 ;
        RECT 52.875 141.375 53.115 141.450 ;
        RECT 50.985 141.055 52.350 141.225 ;
        RECT 50.985 140.655 51.245 141.055 ;
      LAYER mcon ;
        RECT 32.915 173.515 33.085 173.685 ;
        RECT 38.065 172.915 38.235 173.085 ;
        RECT 38.515 170.665 38.685 170.835 ;
        RECT 40.615 170.665 40.785 170.835 ;
        RECT 29.465 168.365 29.635 168.535 ;
        RECT 52.640 162.500 52.840 162.700 ;
        RECT 50.115 162.075 50.285 162.245 ;
        RECT 50.530 162.045 50.700 162.215 ;
        RECT 31.365 159.215 31.535 159.385 ;
        RECT 39.085 157.850 39.285 158.050 ;
        RECT 38.255 157.005 38.445 157.195 ;
        RECT 41.065 157.015 41.235 157.185 ;
        RECT 28.415 154.665 28.585 154.835 ;
        RECT 31.360 154.610 31.540 154.790 ;
        RECT 21.615 143.315 21.785 143.485 ;
        RECT 37.465 143.515 37.635 143.685 ;
        RECT 25.315 143.265 25.485 143.435 ;
        RECT 24.365 142.715 24.535 142.885 ;
        RECT 50.115 141.465 50.285 141.635 ;
        RECT 54.015 141.465 54.185 141.635 ;
      LAYER met1 ;
        RECT 32.885 178.285 37.365 178.515 ;
        RECT 32.885 173.455 33.115 178.285 ;
        RECT 32.335 171.185 36.365 171.415 ;
        RECT 29.405 168.550 29.695 168.565 ;
        RECT 24.450 168.350 29.695 168.550 ;
        RECT 24.450 154.850 24.650 168.350 ;
        RECT 29.405 168.335 29.695 168.350 ;
        RECT 32.335 168.185 32.565 171.185 ;
        RECT 36.135 168.665 36.365 171.185 ;
        RECT 37.135 170.865 37.365 178.285 ;
        RECT 40.050 173.900 44.600 174.100 ;
        RECT 38.005 173.100 38.295 173.115 ;
        RECT 40.050 173.100 40.250 173.900 ;
        RECT 38.000 172.900 40.250 173.100 ;
        RECT 38.005 172.885 38.295 172.900 ;
        RECT 37.135 170.635 38.745 170.865 ;
        RECT 40.585 168.665 40.815 170.895 ;
        RECT 36.135 168.435 40.815 168.665 ;
        RECT 31.335 162.535 37.665 162.765 ;
        RECT 31.335 159.155 31.565 162.535 ;
        RECT 31.335 157.285 35.815 157.515 ;
        RECT 28.355 154.850 28.645 154.865 ;
        RECT 24.450 154.650 28.645 154.850 ;
        RECT 31.335 154.820 31.565 157.285 ;
        RECT 24.450 149.000 24.650 154.650 ;
        RECT 28.355 154.635 28.645 154.650 ;
        RECT 31.330 154.580 31.570 154.820 ;
        RECT 31.335 154.435 31.565 154.580 ;
        RECT 35.585 154.515 35.815 157.285 ;
        RECT 37.435 157.215 37.665 162.535 ;
        RECT 44.400 162.550 44.600 173.900 ;
        RECT 47.200 166.350 60.050 166.550 ;
        RECT 47.200 162.550 47.400 166.350 ;
        RECT 52.550 162.550 54.300 162.750 ;
        RECT 44.400 162.350 49.050 162.550 ;
        RECT 52.580 162.470 52.900 162.550 ;
        RECT 48.775 162.335 49.050 162.350 ;
        RECT 48.775 162.275 50.275 162.335 ;
        RECT 48.775 162.185 50.345 162.275 ;
        RECT 50.055 162.045 50.345 162.185 ;
        RECT 50.500 162.200 50.730 162.275 ;
        RECT 50.500 162.050 51.075 162.200 ;
        RECT 50.500 161.985 50.730 162.050 ;
        RECT 50.500 161.700 50.700 161.985 ;
        RECT 38.250 161.500 50.700 161.700 ;
        RECT 38.250 158.050 38.450 161.500 ;
        RECT 39.055 158.050 39.315 158.080 ;
        RECT 38.250 157.850 39.400 158.050 ;
        RECT 39.055 157.820 39.315 157.850 ;
        RECT 38.195 157.215 38.505 157.225 ;
        RECT 37.435 156.985 38.505 157.215 ;
        RECT 41.005 156.985 41.965 157.215 ;
        RECT 38.195 156.975 38.505 156.985 ;
        RECT 41.735 154.515 41.965 156.985 ;
        RECT 35.585 154.285 41.965 154.515 ;
        RECT 54.100 150.500 54.300 162.550 ;
        RECT 19.100 148.800 24.650 149.000 ;
        RECT 35.850 150.300 54.300 150.500 ;
        RECT 19.100 140.100 19.300 148.800 ;
        RECT 21.600 146.550 34.150 146.750 ;
        RECT 21.600 143.545 21.800 146.550 ;
        RECT 21.585 143.255 21.815 143.545 ;
        RECT 25.255 143.450 25.545 143.465 ;
        RECT 25.255 143.250 26.750 143.450 ;
        RECT 25.255 143.235 25.545 143.250 ;
        RECT 24.305 142.900 24.595 142.915 ;
        RECT 24.305 142.700 25.800 142.900 ;
        RECT 24.305 142.685 24.595 142.700 ;
        RECT 25.600 140.100 25.800 142.700 ;
        RECT 26.550 141.300 26.750 143.250 ;
        RECT 26.550 141.100 31.400 141.300 ;
        RECT 19.100 139.900 25.800 140.100 ;
        RECT 31.200 139.050 31.400 141.100 ;
        RECT 33.950 141.150 34.150 146.550 ;
        RECT 35.850 143.860 36.050 150.300 ;
        RECT 35.820 143.540 36.080 143.860 ;
        RECT 37.405 143.700 37.695 143.715 ;
        RECT 37.405 143.500 39.350 143.700 ;
        RECT 37.405 143.485 37.695 143.500 ;
        RECT 39.150 141.150 39.350 143.500 ;
        RECT 42.650 142.150 42.850 150.300 ;
        RECT 59.850 148.550 60.050 166.350 ;
        RECT 45.400 148.350 60.050 148.550 ;
        RECT 45.400 145.050 45.600 148.350 ;
        RECT 45.400 144.850 54.200 145.050 ;
        RECT 44.320 142.150 44.580 142.210 ;
        RECT 42.650 141.950 44.580 142.150 ;
        RECT 44.320 141.890 44.580 141.950 ;
        RECT 33.950 140.950 39.350 141.150 ;
        RECT 45.400 139.050 45.600 144.850 ;
        RECT 46.420 142.150 46.680 142.210 ;
        RECT 46.420 141.950 50.300 142.150 ;
        RECT 46.420 141.890 46.680 141.950 ;
        RECT 50.100 141.695 50.300 141.950 ;
        RECT 54.000 141.695 54.200 144.850 ;
        RECT 50.085 141.405 50.315 141.695 ;
        RECT 53.985 141.405 54.215 141.695 ;
        RECT 31.200 138.850 45.600 139.050 ;
      LAYER via ;
        RECT 44.320 141.920 44.580 142.180 ;
        RECT 46.420 141.920 46.680 142.180 ;
      LAYER met2 ;
        RECT 44.290 142.150 44.610 142.180 ;
        RECT 46.390 142.150 46.710 142.180 ;
        RECT 44.290 141.950 46.710 142.150 ;
        RECT 44.290 141.920 44.610 141.950 ;
        RECT 46.390 141.920 46.710 141.950 ;
  END
END tt_um_test_8
END LIBRARY

