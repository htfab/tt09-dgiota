VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DIGI_OTA
  CLASS BLOCK ;
  FOREIGN tt_um_DIGI_OTA ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN Out
    ANTENNADIFFAREA 0.601000 ;
    PORT
      LAYER li1 ;
        RECT 53.885 105.895 55.505 106.865 ;
        RECT 53.885 105.225 54.225 105.895 ;
        RECT 53.885 104.655 54.355 105.225 ;
      LAYER mcon ;
        RECT 53.945 105.165 54.115 105.335 ;
      LAYER met1 ;
        RECT 53.870 105.120 54.190 105.380 ;
      LAYER via ;
        RECT 53.900 105.120 54.160 105.380 ;
      LAYER met2 ;
        RECT 53.900 105.090 54.160 105.410 ;
        RECT 53.960 104.925 54.100 105.090 ;
        RECT 53.890 104.555 54.170 104.925 ;
      LAYER via2 ;
        RECT 53.890 104.600 54.170 104.880 ;
      LAYER met3 ;
        RECT 32.160 105.140 33.060 105.190 ;
        RECT 32.160 105.040 33.720 105.140 ;
        RECT 30.230 104.890 42.000 105.040 ;
        RECT 53.865 104.890 54.195 104.905 ;
        RECT 30.230 104.590 54.195 104.890 ;
        RECT 30.230 104.440 42.000 104.590 ;
        RECT 53.865 104.575 54.195 104.590 ;
        RECT 32.160 104.290 33.720 104.440 ;
        RECT 32.820 104.240 33.720 104.290 ;
      LAYER via3 ;
        RECT 32.250 104.380 32.970 105.100 ;
      LAYER met4 ;
        RECT 27.800 161.470 152.710 162.370 ;
        RECT 27.800 105.140 28.700 161.470 ;
        RECT 32.155 105.140 33.065 105.195 ;
        RECT 27.800 104.240 33.720 105.140 ;
        RECT 151.810 0.000 152.710 161.470 ;
    END
  END Out
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN VDPWR
    ANTENNAGATEAREA 1069.782959 ;
    ANTENNADIFFAREA 255.487289 ;
    PORT
      LAYER nwell ;
        RECT 45.330 132.905 134.490 135.735 ;
        RECT 45.330 127.465 134.490 130.295 ;
        RECT 45.330 122.025 134.490 124.855 ;
        RECT 45.330 116.585 134.490 119.415 ;
        RECT 45.330 111.145 134.490 113.975 ;
        RECT 45.330 105.705 134.490 108.535 ;
        RECT 45.330 100.265 134.490 103.095 ;
        RECT 45.330 94.825 134.490 97.655 ;
        RECT 45.330 89.385 134.490 92.215 ;
        RECT 45.330 83.945 134.490 86.775 ;
        RECT 45.330 78.505 134.490 81.335 ;
        RECT 45.330 73.065 134.490 75.895 ;
        RECT 45.330 67.625 134.490 70.455 ;
        RECT 45.330 62.185 134.490 65.015 ;
      LAYER li1 ;
        RECT 46.295 135.495 46.815 136.035 ;
        RECT 45.605 134.405 46.815 135.495 ;
        RECT 50.390 134.840 50.740 136.090 ;
        RECT 55.910 134.840 56.260 136.090 ;
        RECT 46.985 134.405 52.330 134.840 ;
        RECT 52.505 134.405 57.850 134.840 ;
        RECT 58.485 134.405 58.775 135.570 ;
        RECT 62.350 134.840 62.700 136.090 ;
        RECT 67.870 134.840 68.220 136.090 ;
        RECT 70.675 135.495 71.195 136.035 ;
        RECT 58.945 134.405 64.290 134.840 ;
        RECT 64.465 134.405 69.810 134.840 ;
        RECT 69.985 134.405 71.195 135.495 ;
        RECT 71.365 134.405 71.655 135.570 ;
        RECT 75.230 134.840 75.580 136.090 ;
        RECT 80.750 134.840 81.100 136.090 ;
        RECT 83.555 135.495 84.075 136.035 ;
        RECT 71.825 134.405 77.170 134.840 ;
        RECT 77.345 134.405 82.690 134.840 ;
        RECT 82.865 134.405 84.075 135.495 ;
        RECT 84.245 134.405 84.535 135.570 ;
        RECT 88.110 134.840 88.460 136.090 ;
        RECT 93.630 134.840 93.980 136.090 ;
        RECT 96.435 135.495 96.955 136.035 ;
        RECT 84.705 134.405 90.050 134.840 ;
        RECT 90.225 134.405 95.570 134.840 ;
        RECT 95.745 134.405 96.955 135.495 ;
        RECT 97.125 134.405 97.415 135.570 ;
        RECT 100.990 134.840 101.340 136.090 ;
        RECT 106.510 134.840 106.860 136.090 ;
        RECT 109.315 135.495 109.835 136.035 ;
        RECT 97.585 134.405 102.930 134.840 ;
        RECT 103.105 134.405 108.450 134.840 ;
        RECT 108.625 134.405 109.835 135.495 ;
        RECT 110.005 134.405 110.295 135.570 ;
        RECT 113.870 134.840 114.220 136.090 ;
        RECT 119.390 134.840 119.740 136.090 ;
        RECT 122.195 135.495 122.715 136.035 ;
        RECT 110.465 134.405 115.810 134.840 ;
        RECT 115.985 134.405 121.330 134.840 ;
        RECT 121.505 134.405 122.715 135.495 ;
        RECT 122.885 134.405 123.175 135.570 ;
        RECT 126.750 134.840 127.100 136.090 ;
        RECT 130.685 135.495 132.375 136.015 ;
        RECT 123.345 134.405 128.690 134.840 ;
        RECT 128.865 134.405 132.375 135.495 ;
        RECT 133.005 135.495 133.525 136.035 ;
        RECT 133.005 134.405 134.215 135.495 ;
        RECT 45.520 134.235 134.300 134.405 ;
        RECT 45.605 133.145 46.815 134.235 ;
        RECT 46.985 133.800 52.330 134.235 ;
        RECT 52.505 133.800 57.850 134.235 ;
        RECT 46.295 132.605 46.815 133.145 ;
        RECT 50.390 132.550 50.740 133.800 ;
        RECT 55.910 132.550 56.260 133.800 ;
        RECT 58.485 133.070 58.775 134.235 ;
        RECT 58.945 133.800 64.290 134.235 ;
        RECT 64.465 133.800 69.810 134.235 ;
        RECT 69.985 133.800 75.330 134.235 ;
        RECT 75.505 133.800 80.850 134.235 ;
        RECT 62.350 132.550 62.700 133.800 ;
        RECT 67.870 132.550 68.220 133.800 ;
        RECT 73.390 132.550 73.740 133.800 ;
        RECT 78.910 132.550 79.260 133.800 ;
        RECT 81.025 133.145 83.615 134.235 ;
        RECT 82.405 132.625 83.615 133.145 ;
        RECT 84.245 133.070 84.535 134.235 ;
        RECT 84.705 133.800 90.050 134.235 ;
        RECT 90.225 133.800 95.570 134.235 ;
        RECT 95.745 133.800 101.090 134.235 ;
        RECT 101.265 133.800 106.610 134.235 ;
        RECT 88.110 132.550 88.460 133.800 ;
        RECT 93.630 132.550 93.980 133.800 ;
        RECT 99.150 132.550 99.500 133.800 ;
        RECT 104.670 132.550 105.020 133.800 ;
        RECT 106.785 133.145 109.375 134.235 ;
        RECT 108.165 132.625 109.375 133.145 ;
        RECT 110.005 133.070 110.295 134.235 ;
        RECT 110.465 133.800 115.810 134.235 ;
        RECT 115.985 133.800 121.330 134.235 ;
        RECT 121.505 133.800 126.850 134.235 ;
        RECT 127.025 133.800 132.370 134.235 ;
        RECT 113.870 132.550 114.220 133.800 ;
        RECT 119.390 132.550 119.740 133.800 ;
        RECT 124.910 132.550 125.260 133.800 ;
        RECT 130.430 132.550 130.780 133.800 ;
        RECT 133.005 133.145 134.215 134.235 ;
        RECT 133.005 132.605 133.525 133.145 ;
        RECT 46.295 130.055 46.815 130.595 ;
        RECT 45.605 128.965 46.815 130.055 ;
        RECT 50.390 129.400 50.740 130.650 ;
        RECT 55.910 129.400 56.260 130.650 ;
        RECT 61.430 129.400 61.780 130.650 ;
        RECT 66.950 129.400 67.300 130.650 ;
        RECT 69.985 130.055 70.735 130.575 ;
        RECT 46.985 128.965 52.330 129.400 ;
        RECT 52.505 128.965 57.850 129.400 ;
        RECT 58.025 128.965 63.370 129.400 ;
        RECT 63.545 128.965 68.890 129.400 ;
        RECT 69.065 128.965 70.735 130.055 ;
        RECT 71.365 128.965 71.655 130.130 ;
        RECT 75.230 129.400 75.580 130.650 ;
        RECT 80.750 129.400 81.100 130.650 ;
        RECT 86.270 129.400 86.620 130.650 ;
        RECT 91.790 129.400 92.140 130.650 ;
        RECT 95.285 130.055 96.495 130.575 ;
        RECT 71.825 128.965 77.170 129.400 ;
        RECT 77.345 128.965 82.690 129.400 ;
        RECT 82.865 128.965 88.210 129.400 ;
        RECT 88.385 128.965 93.730 129.400 ;
        RECT 93.905 128.965 96.495 130.055 ;
        RECT 97.125 128.965 97.415 130.130 ;
        RECT 100.990 129.400 101.340 130.650 ;
        RECT 106.510 129.400 106.860 130.650 ;
        RECT 112.030 129.400 112.380 130.650 ;
        RECT 117.550 129.400 117.900 130.650 ;
        RECT 121.045 130.055 122.255 130.575 ;
        RECT 97.585 128.965 102.930 129.400 ;
        RECT 103.105 128.965 108.450 129.400 ;
        RECT 108.625 128.965 113.970 129.400 ;
        RECT 114.145 128.965 119.490 129.400 ;
        RECT 119.665 128.965 122.255 130.055 ;
        RECT 122.885 128.965 123.175 130.130 ;
        RECT 126.750 129.400 127.100 130.650 ;
        RECT 130.685 130.055 132.375 130.575 ;
        RECT 123.345 128.965 128.690 129.400 ;
        RECT 128.865 128.965 132.375 130.055 ;
        RECT 133.005 130.055 133.525 130.595 ;
        RECT 133.005 128.965 134.215 130.055 ;
        RECT 45.520 128.795 134.300 128.965 ;
        RECT 45.605 127.705 46.815 128.795 ;
        RECT 46.985 128.360 52.330 128.795 ;
        RECT 52.505 128.360 57.850 128.795 ;
        RECT 46.295 127.165 46.815 127.705 ;
        RECT 50.390 127.110 50.740 128.360 ;
        RECT 55.910 127.110 56.260 128.360 ;
        RECT 58.485 127.630 58.775 128.795 ;
        RECT 58.945 128.360 64.290 128.795 ;
        RECT 64.465 128.360 69.810 128.795 ;
        RECT 69.985 128.360 75.330 128.795 ;
        RECT 75.505 128.360 80.850 128.795 ;
        RECT 62.350 127.110 62.700 128.360 ;
        RECT 67.870 127.110 68.220 128.360 ;
        RECT 73.390 127.110 73.740 128.360 ;
        RECT 78.910 127.110 79.260 128.360 ;
        RECT 81.025 127.705 83.615 128.795 ;
        RECT 82.405 127.185 83.615 127.705 ;
        RECT 84.245 127.630 84.535 128.795 ;
        RECT 84.705 128.360 90.050 128.795 ;
        RECT 90.225 128.360 95.570 128.795 ;
        RECT 95.745 128.360 101.090 128.795 ;
        RECT 101.265 128.360 106.610 128.795 ;
        RECT 88.110 127.110 88.460 128.360 ;
        RECT 93.630 127.110 93.980 128.360 ;
        RECT 99.150 127.110 99.500 128.360 ;
        RECT 104.670 127.110 105.020 128.360 ;
        RECT 106.785 127.705 109.375 128.795 ;
        RECT 108.165 127.185 109.375 127.705 ;
        RECT 110.005 127.630 110.295 128.795 ;
        RECT 110.465 128.360 115.810 128.795 ;
        RECT 115.985 128.360 121.330 128.795 ;
        RECT 121.505 128.360 126.850 128.795 ;
        RECT 127.025 128.360 132.370 128.795 ;
        RECT 113.870 127.110 114.220 128.360 ;
        RECT 119.390 127.110 119.740 128.360 ;
        RECT 124.910 127.110 125.260 128.360 ;
        RECT 130.430 127.110 130.780 128.360 ;
        RECT 133.005 127.705 134.215 128.795 ;
        RECT 133.005 127.165 133.525 127.705 ;
        RECT 46.295 124.615 46.815 125.155 ;
        RECT 45.605 123.525 46.815 124.615 ;
        RECT 50.390 123.960 50.740 125.210 ;
        RECT 55.910 123.960 56.260 125.210 ;
        RECT 61.430 123.960 61.780 125.210 ;
        RECT 66.950 123.960 67.300 125.210 ;
        RECT 69.985 124.615 70.735 125.135 ;
        RECT 46.985 123.525 52.330 123.960 ;
        RECT 52.505 123.525 57.850 123.960 ;
        RECT 58.025 123.525 63.370 123.960 ;
        RECT 63.545 123.525 68.890 123.960 ;
        RECT 69.065 123.525 70.735 124.615 ;
        RECT 71.365 123.525 71.655 124.690 ;
        RECT 75.230 123.960 75.580 125.210 ;
        RECT 80.750 123.960 81.100 125.210 ;
        RECT 86.270 123.960 86.620 125.210 ;
        RECT 91.790 123.960 92.140 125.210 ;
        RECT 95.285 124.615 96.495 125.135 ;
        RECT 71.825 123.525 77.170 123.960 ;
        RECT 77.345 123.525 82.690 123.960 ;
        RECT 82.865 123.525 88.210 123.960 ;
        RECT 88.385 123.525 93.730 123.960 ;
        RECT 93.905 123.525 96.495 124.615 ;
        RECT 97.125 123.525 97.415 124.690 ;
        RECT 100.990 123.960 101.340 125.210 ;
        RECT 106.510 123.960 106.860 125.210 ;
        RECT 112.030 123.960 112.380 125.210 ;
        RECT 117.550 123.960 117.900 125.210 ;
        RECT 121.045 124.615 122.255 125.135 ;
        RECT 97.585 123.525 102.930 123.960 ;
        RECT 103.105 123.525 108.450 123.960 ;
        RECT 108.625 123.525 113.970 123.960 ;
        RECT 114.145 123.525 119.490 123.960 ;
        RECT 119.665 123.525 122.255 124.615 ;
        RECT 122.885 123.525 123.175 124.690 ;
        RECT 126.750 123.960 127.100 125.210 ;
        RECT 130.685 124.615 132.375 125.135 ;
        RECT 123.345 123.525 128.690 123.960 ;
        RECT 128.865 123.525 132.375 124.615 ;
        RECT 133.005 124.615 133.525 125.155 ;
        RECT 133.005 123.525 134.215 124.615 ;
        RECT 45.520 123.355 134.300 123.525 ;
        RECT 45.605 122.265 46.815 123.355 ;
        RECT 46.985 122.920 52.330 123.355 ;
        RECT 52.505 122.920 57.850 123.355 ;
        RECT 46.295 121.725 46.815 122.265 ;
        RECT 50.390 121.670 50.740 122.920 ;
        RECT 55.910 121.670 56.260 122.920 ;
        RECT 58.485 122.190 58.775 123.355 ;
        RECT 58.945 122.920 64.290 123.355 ;
        RECT 64.465 122.920 69.810 123.355 ;
        RECT 69.985 122.920 75.330 123.355 ;
        RECT 75.505 122.920 80.850 123.355 ;
        RECT 62.350 121.670 62.700 122.920 ;
        RECT 67.870 121.670 68.220 122.920 ;
        RECT 73.390 121.670 73.740 122.920 ;
        RECT 78.910 121.670 79.260 122.920 ;
        RECT 81.025 122.265 83.615 123.355 ;
        RECT 82.405 121.745 83.615 122.265 ;
        RECT 84.245 122.190 84.535 123.355 ;
        RECT 84.705 122.920 90.050 123.355 ;
        RECT 90.225 122.920 95.570 123.355 ;
        RECT 95.745 122.920 101.090 123.355 ;
        RECT 101.265 122.920 106.610 123.355 ;
        RECT 88.110 121.670 88.460 122.920 ;
        RECT 93.630 121.670 93.980 122.920 ;
        RECT 99.150 121.670 99.500 122.920 ;
        RECT 104.670 121.670 105.020 122.920 ;
        RECT 106.785 122.265 109.375 123.355 ;
        RECT 108.165 121.745 109.375 122.265 ;
        RECT 110.005 122.190 110.295 123.355 ;
        RECT 110.465 122.920 115.810 123.355 ;
        RECT 115.985 122.920 121.330 123.355 ;
        RECT 121.505 122.920 126.850 123.355 ;
        RECT 127.025 122.920 132.370 123.355 ;
        RECT 113.870 121.670 114.220 122.920 ;
        RECT 119.390 121.670 119.740 122.920 ;
        RECT 124.910 121.670 125.260 122.920 ;
        RECT 130.430 121.670 130.780 122.920 ;
        RECT 133.005 122.265 134.215 123.355 ;
        RECT 133.005 121.725 133.525 122.265 ;
        RECT 46.295 119.175 46.815 119.715 ;
        RECT 45.605 118.085 46.815 119.175 ;
        RECT 50.390 118.520 50.740 119.770 ;
        RECT 55.910 118.520 56.260 119.770 ;
        RECT 61.430 118.520 61.780 119.770 ;
        RECT 66.950 118.520 67.300 119.770 ;
        RECT 69.985 119.175 70.735 119.695 ;
        RECT 46.985 118.085 52.330 118.520 ;
        RECT 52.505 118.085 57.850 118.520 ;
        RECT 58.025 118.085 63.370 118.520 ;
        RECT 63.545 118.085 68.890 118.520 ;
        RECT 69.065 118.085 70.735 119.175 ;
        RECT 71.365 118.085 71.655 119.250 ;
        RECT 75.230 118.520 75.580 119.770 ;
        RECT 80.750 118.520 81.100 119.770 ;
        RECT 86.270 118.520 86.620 119.770 ;
        RECT 91.790 118.520 92.140 119.770 ;
        RECT 95.285 119.175 96.495 119.695 ;
        RECT 71.825 118.085 77.170 118.520 ;
        RECT 77.345 118.085 82.690 118.520 ;
        RECT 82.865 118.085 88.210 118.520 ;
        RECT 88.385 118.085 93.730 118.520 ;
        RECT 93.905 118.085 96.495 119.175 ;
        RECT 97.125 118.085 97.415 119.250 ;
        RECT 100.990 118.520 101.340 119.770 ;
        RECT 106.510 118.520 106.860 119.770 ;
        RECT 112.030 118.520 112.380 119.770 ;
        RECT 117.550 118.520 117.900 119.770 ;
        RECT 121.045 119.175 122.255 119.695 ;
        RECT 97.585 118.085 102.930 118.520 ;
        RECT 103.105 118.085 108.450 118.520 ;
        RECT 108.625 118.085 113.970 118.520 ;
        RECT 114.145 118.085 119.490 118.520 ;
        RECT 119.665 118.085 122.255 119.175 ;
        RECT 122.885 118.085 123.175 119.250 ;
        RECT 126.750 118.520 127.100 119.770 ;
        RECT 130.685 119.175 132.375 119.695 ;
        RECT 123.345 118.085 128.690 118.520 ;
        RECT 128.865 118.085 132.375 119.175 ;
        RECT 133.005 119.175 133.525 119.715 ;
        RECT 133.005 118.085 134.215 119.175 ;
        RECT 45.520 117.915 134.300 118.085 ;
        RECT 45.605 116.825 46.815 117.915 ;
        RECT 46.985 117.480 52.330 117.915 ;
        RECT 52.505 117.480 57.850 117.915 ;
        RECT 46.295 116.285 46.815 116.825 ;
        RECT 50.390 116.230 50.740 117.480 ;
        RECT 55.910 116.230 56.260 117.480 ;
        RECT 58.485 116.750 58.775 117.915 ;
        RECT 58.945 117.480 64.290 117.915 ;
        RECT 64.465 117.480 69.810 117.915 ;
        RECT 69.985 117.480 75.330 117.915 ;
        RECT 75.505 117.480 80.850 117.915 ;
        RECT 62.350 116.230 62.700 117.480 ;
        RECT 67.870 116.230 68.220 117.480 ;
        RECT 73.390 116.230 73.740 117.480 ;
        RECT 78.910 116.230 79.260 117.480 ;
        RECT 81.025 116.825 83.615 117.915 ;
        RECT 82.405 116.305 83.615 116.825 ;
        RECT 84.245 116.750 84.535 117.915 ;
        RECT 84.705 117.480 90.050 117.915 ;
        RECT 90.225 117.480 95.570 117.915 ;
        RECT 95.745 117.480 101.090 117.915 ;
        RECT 101.265 117.480 106.610 117.915 ;
        RECT 88.110 116.230 88.460 117.480 ;
        RECT 93.630 116.230 93.980 117.480 ;
        RECT 99.150 116.230 99.500 117.480 ;
        RECT 104.670 116.230 105.020 117.480 ;
        RECT 106.785 116.825 109.375 117.915 ;
        RECT 108.165 116.305 109.375 116.825 ;
        RECT 110.005 116.750 110.295 117.915 ;
        RECT 110.465 117.480 115.810 117.915 ;
        RECT 115.985 117.480 121.330 117.915 ;
        RECT 121.505 117.480 126.850 117.915 ;
        RECT 127.025 117.480 132.370 117.915 ;
        RECT 113.870 116.230 114.220 117.480 ;
        RECT 119.390 116.230 119.740 117.480 ;
        RECT 124.910 116.230 125.260 117.480 ;
        RECT 130.430 116.230 130.780 117.480 ;
        RECT 133.005 116.825 134.215 117.915 ;
        RECT 133.005 116.285 133.525 116.825 ;
        RECT 46.295 113.735 46.815 114.275 ;
        RECT 45.605 112.645 46.815 113.735 ;
        RECT 50.390 113.080 50.740 114.330 ;
        RECT 55.910 113.080 56.260 114.330 ;
        RECT 61.430 113.080 61.780 114.330 ;
        RECT 66.950 113.080 67.300 114.330 ;
        RECT 69.985 113.735 70.735 114.255 ;
        RECT 46.985 112.645 52.330 113.080 ;
        RECT 52.505 112.645 57.850 113.080 ;
        RECT 58.025 112.645 63.370 113.080 ;
        RECT 63.545 112.645 68.890 113.080 ;
        RECT 69.065 112.645 70.735 113.735 ;
        RECT 71.365 112.645 71.655 113.810 ;
        RECT 75.230 113.080 75.580 114.330 ;
        RECT 80.750 113.080 81.100 114.330 ;
        RECT 86.270 113.080 86.620 114.330 ;
        RECT 91.790 113.080 92.140 114.330 ;
        RECT 95.285 113.735 96.495 114.255 ;
        RECT 71.825 112.645 77.170 113.080 ;
        RECT 77.345 112.645 82.690 113.080 ;
        RECT 82.865 112.645 88.210 113.080 ;
        RECT 88.385 112.645 93.730 113.080 ;
        RECT 93.905 112.645 96.495 113.735 ;
        RECT 97.125 112.645 97.415 113.810 ;
        RECT 100.990 113.080 101.340 114.330 ;
        RECT 106.510 113.080 106.860 114.330 ;
        RECT 112.030 113.080 112.380 114.330 ;
        RECT 117.550 113.080 117.900 114.330 ;
        RECT 121.045 113.735 122.255 114.255 ;
        RECT 97.585 112.645 102.930 113.080 ;
        RECT 103.105 112.645 108.450 113.080 ;
        RECT 108.625 112.645 113.970 113.080 ;
        RECT 114.145 112.645 119.490 113.080 ;
        RECT 119.665 112.645 122.255 113.735 ;
        RECT 122.885 112.645 123.175 113.810 ;
        RECT 126.750 113.080 127.100 114.330 ;
        RECT 130.685 113.735 132.375 114.255 ;
        RECT 123.345 112.645 128.690 113.080 ;
        RECT 128.865 112.645 132.375 113.735 ;
        RECT 133.005 113.735 133.525 114.275 ;
        RECT 133.005 112.645 134.215 113.735 ;
        RECT 45.520 112.475 134.300 112.645 ;
        RECT 45.605 111.385 46.815 112.475 ;
        RECT 46.985 112.040 52.330 112.475 ;
        RECT 52.505 112.040 57.850 112.475 ;
        RECT 46.295 110.845 46.815 111.385 ;
        RECT 50.390 110.790 50.740 112.040 ;
        RECT 55.910 110.790 56.260 112.040 ;
        RECT 58.485 111.310 58.775 112.475 ;
        RECT 58.945 112.040 64.290 112.475 ;
        RECT 64.465 112.040 69.810 112.475 ;
        RECT 69.985 112.040 75.330 112.475 ;
        RECT 75.505 112.040 80.850 112.475 ;
        RECT 62.350 110.790 62.700 112.040 ;
        RECT 67.870 110.790 68.220 112.040 ;
        RECT 73.390 110.790 73.740 112.040 ;
        RECT 78.910 110.790 79.260 112.040 ;
        RECT 81.025 111.385 83.615 112.475 ;
        RECT 82.405 110.865 83.615 111.385 ;
        RECT 84.245 111.310 84.535 112.475 ;
        RECT 84.705 112.040 90.050 112.475 ;
        RECT 90.225 112.040 95.570 112.475 ;
        RECT 95.745 112.040 101.090 112.475 ;
        RECT 101.265 112.040 106.610 112.475 ;
        RECT 88.110 110.790 88.460 112.040 ;
        RECT 93.630 110.790 93.980 112.040 ;
        RECT 99.150 110.790 99.500 112.040 ;
        RECT 104.670 110.790 105.020 112.040 ;
        RECT 106.785 111.385 109.375 112.475 ;
        RECT 108.165 110.865 109.375 111.385 ;
        RECT 110.005 111.310 110.295 112.475 ;
        RECT 110.465 112.040 115.810 112.475 ;
        RECT 115.985 112.040 121.330 112.475 ;
        RECT 121.505 112.040 126.850 112.475 ;
        RECT 127.025 112.040 132.370 112.475 ;
        RECT 113.870 110.790 114.220 112.040 ;
        RECT 119.390 110.790 119.740 112.040 ;
        RECT 124.910 110.790 125.260 112.040 ;
        RECT 130.430 110.790 130.780 112.040 ;
        RECT 133.005 111.385 134.215 112.475 ;
        RECT 133.005 110.845 133.525 111.385 ;
        RECT 46.295 108.295 46.815 108.835 ;
        RECT 45.605 107.205 46.815 108.295 ;
        RECT 50.390 107.640 50.740 108.890 ;
        RECT 55.910 107.640 56.260 108.890 ;
        RECT 58.945 108.295 59.695 108.815 ;
        RECT 46.985 107.205 52.330 107.640 ;
        RECT 52.505 107.205 57.850 107.640 ;
        RECT 58.025 107.205 59.695 108.295 ;
        RECT 60.365 107.205 60.595 108.345 ;
        RECT 61.265 107.205 61.475 108.345 ;
        RECT 62.180 107.205 62.510 107.965 ;
        RECT 63.110 107.205 63.370 108.355 ;
        RECT 66.950 107.640 67.300 108.890 ;
        RECT 69.985 108.295 70.735 108.815 ;
        RECT 63.545 107.205 68.890 107.640 ;
        RECT 69.065 107.205 70.735 108.295 ;
        RECT 71.365 107.205 71.655 108.370 ;
        RECT 75.230 107.640 75.580 108.890 ;
        RECT 80.750 107.640 81.100 108.890 ;
        RECT 86.270 107.640 86.620 108.890 ;
        RECT 91.790 107.640 92.140 108.890 ;
        RECT 95.285 108.295 96.495 108.815 ;
        RECT 71.825 107.205 77.170 107.640 ;
        RECT 77.345 107.205 82.690 107.640 ;
        RECT 82.865 107.205 88.210 107.640 ;
        RECT 88.385 107.205 93.730 107.640 ;
        RECT 93.905 107.205 96.495 108.295 ;
        RECT 97.125 107.205 97.415 108.370 ;
        RECT 100.990 107.640 101.340 108.890 ;
        RECT 106.510 107.640 106.860 108.890 ;
        RECT 112.030 107.640 112.380 108.890 ;
        RECT 117.550 107.640 117.900 108.890 ;
        RECT 121.045 108.295 122.255 108.815 ;
        RECT 97.585 107.205 102.930 107.640 ;
        RECT 103.105 107.205 108.450 107.640 ;
        RECT 108.625 107.205 113.970 107.640 ;
        RECT 114.145 107.205 119.490 107.640 ;
        RECT 119.665 107.205 122.255 108.295 ;
        RECT 122.885 107.205 123.175 108.370 ;
        RECT 126.750 107.640 127.100 108.890 ;
        RECT 130.685 108.295 132.375 108.815 ;
        RECT 123.345 107.205 128.690 107.640 ;
        RECT 128.865 107.205 132.375 108.295 ;
        RECT 133.005 108.295 133.525 108.835 ;
        RECT 133.005 107.205 134.215 108.295 ;
        RECT 45.520 107.035 134.300 107.205 ;
        RECT 45.605 105.945 46.815 107.035 ;
        RECT 46.985 105.945 50.495 107.035 ;
        RECT 46.295 105.405 46.815 105.945 ;
        RECT 48.805 105.425 50.495 105.945 ;
        RECT 51.185 105.895 51.395 107.035 ;
        RECT 52.065 105.895 52.295 107.035 ;
        RECT 52.505 105.895 52.785 107.035 ;
        RECT 53.455 105.895 53.715 107.035 ;
        RECT 55.675 106.575 56.040 107.035 ;
        RECT 56.635 106.575 56.965 107.035 ;
        RECT 58.485 105.870 58.775 107.035 ;
        RECT 58.945 106.600 64.290 107.035 ;
        RECT 64.465 106.600 69.810 107.035 ;
        RECT 69.985 106.600 75.330 107.035 ;
        RECT 75.505 106.600 80.850 107.035 ;
        RECT 62.350 105.350 62.700 106.600 ;
        RECT 67.870 105.350 68.220 106.600 ;
        RECT 73.390 105.350 73.740 106.600 ;
        RECT 78.910 105.350 79.260 106.600 ;
        RECT 81.025 105.945 83.615 107.035 ;
        RECT 82.405 105.425 83.615 105.945 ;
        RECT 84.245 105.870 84.535 107.035 ;
        RECT 84.705 106.600 90.050 107.035 ;
        RECT 90.225 106.600 95.570 107.035 ;
        RECT 95.745 106.600 101.090 107.035 ;
        RECT 101.265 106.600 106.610 107.035 ;
        RECT 88.110 105.350 88.460 106.600 ;
        RECT 93.630 105.350 93.980 106.600 ;
        RECT 99.150 105.350 99.500 106.600 ;
        RECT 104.670 105.350 105.020 106.600 ;
        RECT 106.785 105.945 109.375 107.035 ;
        RECT 108.165 105.425 109.375 105.945 ;
        RECT 110.005 105.870 110.295 107.035 ;
        RECT 110.465 106.600 115.810 107.035 ;
        RECT 115.985 106.600 121.330 107.035 ;
        RECT 121.505 106.600 126.850 107.035 ;
        RECT 127.025 106.600 132.370 107.035 ;
        RECT 113.870 105.350 114.220 106.600 ;
        RECT 119.390 105.350 119.740 106.600 ;
        RECT 124.910 105.350 125.260 106.600 ;
        RECT 130.430 105.350 130.780 106.600 ;
        RECT 133.005 105.945 134.215 107.035 ;
        RECT 133.005 105.405 133.525 105.945 ;
        RECT 46.295 102.855 46.815 103.395 ;
        RECT 45.605 101.765 46.815 102.855 ;
        RECT 47.425 101.765 47.755 102.525 ;
        RECT 51.770 102.200 52.120 103.450 ;
        RECT 48.365 101.765 53.710 102.200 ;
        RECT 54.805 101.765 55.065 102.905 ;
        RECT 55.735 101.765 55.905 102.565 ;
        RECT 56.575 101.765 56.830 102.565 ;
        RECT 57.535 101.765 57.970 102.555 ;
        RECT 64.650 102.200 65.000 103.450 ;
        RECT 68.585 102.855 70.275 103.375 ;
        RECT 59.000 101.765 59.330 102.125 ;
        RECT 61.245 101.765 66.590 102.200 ;
        RECT 66.765 101.765 70.275 102.855 ;
        RECT 71.365 101.765 71.655 102.930 ;
        RECT 75.230 102.200 75.580 103.450 ;
        RECT 80.750 102.200 81.100 103.450 ;
        RECT 86.270 102.200 86.620 103.450 ;
        RECT 91.790 102.200 92.140 103.450 ;
        RECT 95.285 102.855 96.495 103.375 ;
        RECT 71.825 101.765 77.170 102.200 ;
        RECT 77.345 101.765 82.690 102.200 ;
        RECT 82.865 101.765 88.210 102.200 ;
        RECT 88.385 101.765 93.730 102.200 ;
        RECT 93.905 101.765 96.495 102.855 ;
        RECT 97.125 101.765 97.415 102.930 ;
        RECT 100.990 102.200 101.340 103.450 ;
        RECT 106.510 102.200 106.860 103.450 ;
        RECT 112.030 102.200 112.380 103.450 ;
        RECT 117.550 102.200 117.900 103.450 ;
        RECT 121.045 102.855 122.255 103.375 ;
        RECT 97.585 101.765 102.930 102.200 ;
        RECT 103.105 101.765 108.450 102.200 ;
        RECT 108.625 101.765 113.970 102.200 ;
        RECT 114.145 101.765 119.490 102.200 ;
        RECT 119.665 101.765 122.255 102.855 ;
        RECT 122.885 101.765 123.175 102.930 ;
        RECT 126.750 102.200 127.100 103.450 ;
        RECT 130.685 102.855 132.375 103.375 ;
        RECT 123.345 101.765 128.690 102.200 ;
        RECT 128.865 101.765 132.375 102.855 ;
        RECT 133.005 102.855 133.525 103.395 ;
        RECT 133.005 101.765 134.215 102.855 ;
        RECT 45.520 101.595 134.300 101.765 ;
        RECT 45.605 100.505 46.815 101.595 ;
        RECT 47.425 100.835 47.755 101.595 ;
        RECT 48.365 101.160 53.710 101.595 ;
        RECT 46.295 99.965 46.815 100.505 ;
        RECT 51.770 99.910 52.120 101.160 ;
        RECT 53.885 100.505 57.395 101.595 ;
        RECT 55.705 99.985 57.395 100.505 ;
        RECT 58.485 100.430 58.775 101.595 ;
        RECT 58.945 101.160 64.290 101.595 ;
        RECT 64.465 101.160 69.810 101.595 ;
        RECT 69.985 101.160 75.330 101.595 ;
        RECT 75.505 101.160 80.850 101.595 ;
        RECT 62.350 99.910 62.700 101.160 ;
        RECT 67.870 99.910 68.220 101.160 ;
        RECT 73.390 99.910 73.740 101.160 ;
        RECT 78.910 99.910 79.260 101.160 ;
        RECT 81.025 100.505 83.615 101.595 ;
        RECT 82.405 99.985 83.615 100.505 ;
        RECT 84.245 100.430 84.535 101.595 ;
        RECT 84.705 101.160 90.050 101.595 ;
        RECT 90.225 101.160 95.570 101.595 ;
        RECT 95.745 101.160 101.090 101.595 ;
        RECT 101.265 101.160 106.610 101.595 ;
        RECT 88.110 99.910 88.460 101.160 ;
        RECT 93.630 99.910 93.980 101.160 ;
        RECT 99.150 99.910 99.500 101.160 ;
        RECT 104.670 99.910 105.020 101.160 ;
        RECT 106.785 100.505 109.375 101.595 ;
        RECT 108.165 99.985 109.375 100.505 ;
        RECT 110.005 100.430 110.295 101.595 ;
        RECT 110.465 101.160 115.810 101.595 ;
        RECT 115.985 101.160 121.330 101.595 ;
        RECT 121.505 101.160 126.850 101.595 ;
        RECT 127.025 101.160 132.370 101.595 ;
        RECT 113.870 99.910 114.220 101.160 ;
        RECT 119.390 99.910 119.740 101.160 ;
        RECT 124.910 99.910 125.260 101.160 ;
        RECT 130.430 99.910 130.780 101.160 ;
        RECT 133.005 100.505 134.215 101.595 ;
        RECT 133.005 99.965 133.525 100.505 ;
        RECT 46.295 97.415 46.815 97.955 ;
        RECT 45.605 96.325 46.815 97.415 ;
        RECT 50.390 96.760 50.740 98.010 ;
        RECT 53.885 97.415 55.095 97.935 ;
        RECT 46.985 96.325 52.330 96.760 ;
        RECT 52.505 96.325 55.095 97.415 ;
        RECT 56.165 96.325 56.495 97.085 ;
        RECT 60.510 96.760 60.860 98.010 ;
        RECT 66.030 96.760 66.380 98.010 ;
        RECT 69.525 97.415 70.735 97.935 ;
        RECT 57.105 96.325 62.450 96.760 ;
        RECT 62.625 96.325 67.970 96.760 ;
        RECT 68.145 96.325 70.735 97.415 ;
        RECT 71.365 96.325 71.655 97.490 ;
        RECT 75.230 96.760 75.580 98.010 ;
        RECT 80.750 96.760 81.100 98.010 ;
        RECT 86.270 96.760 86.620 98.010 ;
        RECT 91.790 96.760 92.140 98.010 ;
        RECT 95.285 97.415 96.495 97.935 ;
        RECT 71.825 96.325 77.170 96.760 ;
        RECT 77.345 96.325 82.690 96.760 ;
        RECT 82.865 96.325 88.210 96.760 ;
        RECT 88.385 96.325 93.730 96.760 ;
        RECT 93.905 96.325 96.495 97.415 ;
        RECT 97.125 96.325 97.415 97.490 ;
        RECT 100.990 96.760 101.340 98.010 ;
        RECT 106.510 96.760 106.860 98.010 ;
        RECT 112.030 96.760 112.380 98.010 ;
        RECT 117.550 96.760 117.900 98.010 ;
        RECT 121.045 97.415 122.255 97.935 ;
        RECT 97.585 96.325 102.930 96.760 ;
        RECT 103.105 96.325 108.450 96.760 ;
        RECT 108.625 96.325 113.970 96.760 ;
        RECT 114.145 96.325 119.490 96.760 ;
        RECT 119.665 96.325 122.255 97.415 ;
        RECT 122.885 96.325 123.175 97.490 ;
        RECT 126.750 96.760 127.100 98.010 ;
        RECT 130.685 97.415 132.375 97.935 ;
        RECT 123.345 96.325 128.690 96.760 ;
        RECT 128.865 96.325 132.375 97.415 ;
        RECT 133.005 97.415 133.525 97.955 ;
        RECT 133.005 96.325 134.215 97.415 ;
        RECT 45.520 96.155 134.300 96.325 ;
        RECT 45.605 95.065 46.815 96.155 ;
        RECT 46.985 95.720 52.330 96.155 ;
        RECT 46.295 94.525 46.815 95.065 ;
        RECT 50.390 94.470 50.740 95.720 ;
        RECT 52.505 95.065 56.015 96.155 ;
        RECT 54.325 94.545 56.015 95.065 ;
        RECT 56.645 95.015 56.905 96.155 ;
        RECT 57.575 95.015 57.855 96.155 ;
        RECT 58.485 94.990 58.775 96.155 ;
        RECT 58.945 95.720 64.290 96.155 ;
        RECT 64.465 95.720 69.810 96.155 ;
        RECT 69.985 95.720 75.330 96.155 ;
        RECT 75.505 95.720 80.850 96.155 ;
        RECT 62.350 94.470 62.700 95.720 ;
        RECT 67.870 94.470 68.220 95.720 ;
        RECT 73.390 94.470 73.740 95.720 ;
        RECT 78.910 94.470 79.260 95.720 ;
        RECT 81.025 95.065 83.615 96.155 ;
        RECT 82.405 94.545 83.615 95.065 ;
        RECT 84.245 94.990 84.535 96.155 ;
        RECT 84.705 95.720 90.050 96.155 ;
        RECT 90.225 95.720 95.570 96.155 ;
        RECT 95.745 95.720 101.090 96.155 ;
        RECT 101.265 95.720 106.610 96.155 ;
        RECT 88.110 94.470 88.460 95.720 ;
        RECT 93.630 94.470 93.980 95.720 ;
        RECT 99.150 94.470 99.500 95.720 ;
        RECT 104.670 94.470 105.020 95.720 ;
        RECT 106.785 95.065 109.375 96.155 ;
        RECT 108.165 94.545 109.375 95.065 ;
        RECT 110.005 94.990 110.295 96.155 ;
        RECT 110.465 95.720 115.810 96.155 ;
        RECT 115.985 95.720 121.330 96.155 ;
        RECT 121.505 95.720 126.850 96.155 ;
        RECT 127.025 95.720 132.370 96.155 ;
        RECT 113.870 94.470 114.220 95.720 ;
        RECT 119.390 94.470 119.740 95.720 ;
        RECT 124.910 94.470 125.260 95.720 ;
        RECT 130.430 94.470 130.780 95.720 ;
        RECT 133.005 95.065 134.215 96.155 ;
        RECT 133.005 94.525 133.525 95.065 ;
        RECT 46.295 91.975 46.815 92.515 ;
        RECT 48.805 91.975 50.495 92.495 ;
        RECT 45.605 90.885 46.815 91.975 ;
        RECT 46.985 90.885 50.495 91.975 ;
        RECT 52.335 90.885 52.505 91.645 ;
        RECT 54.875 90.885 55.045 92.025 ;
        RECT 56.235 90.885 56.405 92.025 ;
        RECT 58.775 90.885 58.945 91.645 ;
        RECT 59.905 90.885 60.135 92.025 ;
        RECT 60.805 90.885 61.015 92.025 ;
        RECT 61.285 90.885 61.515 92.025 ;
        RECT 62.185 90.885 62.395 92.025 ;
        RECT 66.030 91.320 66.380 92.570 ;
        RECT 69.525 91.975 70.735 92.495 ;
        RECT 62.625 90.885 67.970 91.320 ;
        RECT 68.145 90.885 70.735 91.975 ;
        RECT 71.365 90.885 71.655 92.050 ;
        RECT 75.230 91.320 75.580 92.570 ;
        RECT 80.750 91.320 81.100 92.570 ;
        RECT 86.270 91.320 86.620 92.570 ;
        RECT 91.790 91.320 92.140 92.570 ;
        RECT 95.285 91.975 96.495 92.495 ;
        RECT 71.825 90.885 77.170 91.320 ;
        RECT 77.345 90.885 82.690 91.320 ;
        RECT 82.865 90.885 88.210 91.320 ;
        RECT 88.385 90.885 93.730 91.320 ;
        RECT 93.905 90.885 96.495 91.975 ;
        RECT 97.125 90.885 97.415 92.050 ;
        RECT 100.990 91.320 101.340 92.570 ;
        RECT 106.510 91.320 106.860 92.570 ;
        RECT 112.030 91.320 112.380 92.570 ;
        RECT 117.550 91.320 117.900 92.570 ;
        RECT 121.045 91.975 122.255 92.495 ;
        RECT 97.585 90.885 102.930 91.320 ;
        RECT 103.105 90.885 108.450 91.320 ;
        RECT 108.625 90.885 113.970 91.320 ;
        RECT 114.145 90.885 119.490 91.320 ;
        RECT 119.665 90.885 122.255 91.975 ;
        RECT 122.885 90.885 123.175 92.050 ;
        RECT 126.750 91.320 127.100 92.570 ;
        RECT 130.685 91.975 132.375 92.495 ;
        RECT 123.345 90.885 128.690 91.320 ;
        RECT 128.865 90.885 132.375 91.975 ;
        RECT 133.005 91.975 133.525 92.515 ;
        RECT 133.005 90.885 134.215 91.975 ;
        RECT 45.520 90.715 134.300 90.885 ;
        RECT 45.605 89.625 46.815 90.715 ;
        RECT 46.985 90.280 52.330 90.715 ;
        RECT 46.295 89.085 46.815 89.625 ;
        RECT 50.390 89.030 50.740 90.280 ;
        RECT 52.505 89.625 55.095 90.715 ;
        RECT 55.705 89.955 56.035 90.715 ;
        RECT 53.885 89.105 55.095 89.625 ;
        RECT 56.685 89.575 56.915 90.715 ;
        RECT 57.585 89.575 57.795 90.715 ;
        RECT 58.485 89.550 58.775 90.715 ;
        RECT 58.945 90.280 64.290 90.715 ;
        RECT 64.465 90.280 69.810 90.715 ;
        RECT 69.985 90.280 75.330 90.715 ;
        RECT 75.505 90.280 80.850 90.715 ;
        RECT 62.350 89.030 62.700 90.280 ;
        RECT 67.870 89.030 68.220 90.280 ;
        RECT 73.390 89.030 73.740 90.280 ;
        RECT 78.910 89.030 79.260 90.280 ;
        RECT 81.025 89.625 83.615 90.715 ;
        RECT 82.405 89.105 83.615 89.625 ;
        RECT 84.245 89.550 84.535 90.715 ;
        RECT 84.705 90.280 90.050 90.715 ;
        RECT 90.225 90.280 95.570 90.715 ;
        RECT 95.745 90.280 101.090 90.715 ;
        RECT 101.265 90.280 106.610 90.715 ;
        RECT 88.110 89.030 88.460 90.280 ;
        RECT 93.630 89.030 93.980 90.280 ;
        RECT 99.150 89.030 99.500 90.280 ;
        RECT 104.670 89.030 105.020 90.280 ;
        RECT 106.785 89.625 109.375 90.715 ;
        RECT 108.165 89.105 109.375 89.625 ;
        RECT 110.005 89.550 110.295 90.715 ;
        RECT 110.465 90.280 115.810 90.715 ;
        RECT 115.985 90.280 121.330 90.715 ;
        RECT 121.505 90.280 126.850 90.715 ;
        RECT 127.025 90.280 132.370 90.715 ;
        RECT 113.870 89.030 114.220 90.280 ;
        RECT 119.390 89.030 119.740 90.280 ;
        RECT 124.910 89.030 125.260 90.280 ;
        RECT 130.430 89.030 130.780 90.280 ;
        RECT 133.005 89.625 134.215 90.715 ;
        RECT 133.005 89.085 133.525 89.625 ;
        RECT 46.295 86.535 46.815 87.075 ;
        RECT 45.605 85.445 46.815 86.535 ;
        RECT 50.390 85.880 50.740 87.130 ;
        RECT 55.910 85.880 56.260 87.130 ;
        RECT 61.430 85.880 61.780 87.130 ;
        RECT 66.950 85.880 67.300 87.130 ;
        RECT 69.985 86.535 70.735 87.055 ;
        RECT 46.985 85.445 52.330 85.880 ;
        RECT 52.505 85.445 57.850 85.880 ;
        RECT 58.025 85.445 63.370 85.880 ;
        RECT 63.545 85.445 68.890 85.880 ;
        RECT 69.065 85.445 70.735 86.535 ;
        RECT 71.365 85.445 71.655 86.610 ;
        RECT 75.230 85.880 75.580 87.130 ;
        RECT 80.750 85.880 81.100 87.130 ;
        RECT 86.270 85.880 86.620 87.130 ;
        RECT 91.790 85.880 92.140 87.130 ;
        RECT 95.285 86.535 96.495 87.055 ;
        RECT 71.825 85.445 77.170 85.880 ;
        RECT 77.345 85.445 82.690 85.880 ;
        RECT 82.865 85.445 88.210 85.880 ;
        RECT 88.385 85.445 93.730 85.880 ;
        RECT 93.905 85.445 96.495 86.535 ;
        RECT 97.125 85.445 97.415 86.610 ;
        RECT 100.990 85.880 101.340 87.130 ;
        RECT 106.510 85.880 106.860 87.130 ;
        RECT 112.030 85.880 112.380 87.130 ;
        RECT 117.550 85.880 117.900 87.130 ;
        RECT 121.045 86.535 122.255 87.055 ;
        RECT 97.585 85.445 102.930 85.880 ;
        RECT 103.105 85.445 108.450 85.880 ;
        RECT 108.625 85.445 113.970 85.880 ;
        RECT 114.145 85.445 119.490 85.880 ;
        RECT 119.665 85.445 122.255 86.535 ;
        RECT 122.885 85.445 123.175 86.610 ;
        RECT 126.750 85.880 127.100 87.130 ;
        RECT 130.685 86.535 132.375 87.055 ;
        RECT 123.345 85.445 128.690 85.880 ;
        RECT 128.865 85.445 132.375 86.535 ;
        RECT 133.005 86.535 133.525 87.075 ;
        RECT 133.005 85.445 134.215 86.535 ;
        RECT 45.520 85.275 134.300 85.445 ;
        RECT 45.605 84.185 46.815 85.275 ;
        RECT 46.985 84.840 52.330 85.275 ;
        RECT 52.505 84.840 57.850 85.275 ;
        RECT 46.295 83.645 46.815 84.185 ;
        RECT 50.390 83.590 50.740 84.840 ;
        RECT 55.910 83.590 56.260 84.840 ;
        RECT 58.485 84.110 58.775 85.275 ;
        RECT 58.945 84.840 64.290 85.275 ;
        RECT 64.465 84.840 69.810 85.275 ;
        RECT 69.985 84.840 75.330 85.275 ;
        RECT 75.505 84.840 80.850 85.275 ;
        RECT 62.350 83.590 62.700 84.840 ;
        RECT 67.870 83.590 68.220 84.840 ;
        RECT 73.390 83.590 73.740 84.840 ;
        RECT 78.910 83.590 79.260 84.840 ;
        RECT 81.025 84.185 83.615 85.275 ;
        RECT 82.405 83.665 83.615 84.185 ;
        RECT 84.245 84.110 84.535 85.275 ;
        RECT 84.705 84.840 90.050 85.275 ;
        RECT 90.225 84.840 95.570 85.275 ;
        RECT 95.745 84.840 101.090 85.275 ;
        RECT 101.265 84.840 106.610 85.275 ;
        RECT 88.110 83.590 88.460 84.840 ;
        RECT 93.630 83.590 93.980 84.840 ;
        RECT 99.150 83.590 99.500 84.840 ;
        RECT 104.670 83.590 105.020 84.840 ;
        RECT 106.785 84.185 109.375 85.275 ;
        RECT 108.165 83.665 109.375 84.185 ;
        RECT 110.005 84.110 110.295 85.275 ;
        RECT 110.465 84.840 115.810 85.275 ;
        RECT 115.985 84.840 121.330 85.275 ;
        RECT 121.505 84.840 126.850 85.275 ;
        RECT 127.025 84.840 132.370 85.275 ;
        RECT 113.870 83.590 114.220 84.840 ;
        RECT 119.390 83.590 119.740 84.840 ;
        RECT 124.910 83.590 125.260 84.840 ;
        RECT 130.430 83.590 130.780 84.840 ;
        RECT 133.005 84.185 134.215 85.275 ;
        RECT 133.005 83.645 133.525 84.185 ;
        RECT 46.295 81.095 46.815 81.635 ;
        RECT 45.605 80.005 46.815 81.095 ;
        RECT 50.390 80.440 50.740 81.690 ;
        RECT 55.910 80.440 56.260 81.690 ;
        RECT 61.430 80.440 61.780 81.690 ;
        RECT 66.950 80.440 67.300 81.690 ;
        RECT 69.985 81.095 70.735 81.615 ;
        RECT 46.985 80.005 52.330 80.440 ;
        RECT 52.505 80.005 57.850 80.440 ;
        RECT 58.025 80.005 63.370 80.440 ;
        RECT 63.545 80.005 68.890 80.440 ;
        RECT 69.065 80.005 70.735 81.095 ;
        RECT 71.365 80.005 71.655 81.170 ;
        RECT 75.230 80.440 75.580 81.690 ;
        RECT 80.750 80.440 81.100 81.690 ;
        RECT 86.270 80.440 86.620 81.690 ;
        RECT 91.790 80.440 92.140 81.690 ;
        RECT 95.285 81.095 96.495 81.615 ;
        RECT 71.825 80.005 77.170 80.440 ;
        RECT 77.345 80.005 82.690 80.440 ;
        RECT 82.865 80.005 88.210 80.440 ;
        RECT 88.385 80.005 93.730 80.440 ;
        RECT 93.905 80.005 96.495 81.095 ;
        RECT 97.125 80.005 97.415 81.170 ;
        RECT 100.990 80.440 101.340 81.690 ;
        RECT 106.510 80.440 106.860 81.690 ;
        RECT 112.030 80.440 112.380 81.690 ;
        RECT 117.550 80.440 117.900 81.690 ;
        RECT 121.045 81.095 122.255 81.615 ;
        RECT 97.585 80.005 102.930 80.440 ;
        RECT 103.105 80.005 108.450 80.440 ;
        RECT 108.625 80.005 113.970 80.440 ;
        RECT 114.145 80.005 119.490 80.440 ;
        RECT 119.665 80.005 122.255 81.095 ;
        RECT 122.885 80.005 123.175 81.170 ;
        RECT 126.750 80.440 127.100 81.690 ;
        RECT 130.685 81.095 132.375 81.615 ;
        RECT 123.345 80.005 128.690 80.440 ;
        RECT 128.865 80.005 132.375 81.095 ;
        RECT 133.005 81.095 133.525 81.635 ;
        RECT 133.005 80.005 134.215 81.095 ;
        RECT 45.520 79.835 134.300 80.005 ;
        RECT 45.605 78.745 46.815 79.835 ;
        RECT 46.985 79.400 52.330 79.835 ;
        RECT 52.505 79.400 57.850 79.835 ;
        RECT 46.295 78.205 46.815 78.745 ;
        RECT 50.390 78.150 50.740 79.400 ;
        RECT 55.910 78.150 56.260 79.400 ;
        RECT 58.485 78.670 58.775 79.835 ;
        RECT 58.945 79.400 64.290 79.835 ;
        RECT 64.465 79.400 69.810 79.835 ;
        RECT 69.985 79.400 75.330 79.835 ;
        RECT 75.505 79.400 80.850 79.835 ;
        RECT 62.350 78.150 62.700 79.400 ;
        RECT 67.870 78.150 68.220 79.400 ;
        RECT 73.390 78.150 73.740 79.400 ;
        RECT 78.910 78.150 79.260 79.400 ;
        RECT 81.025 78.745 83.615 79.835 ;
        RECT 82.405 78.225 83.615 78.745 ;
        RECT 84.245 78.670 84.535 79.835 ;
        RECT 84.705 79.400 90.050 79.835 ;
        RECT 90.225 79.400 95.570 79.835 ;
        RECT 95.745 79.400 101.090 79.835 ;
        RECT 101.265 79.400 106.610 79.835 ;
        RECT 88.110 78.150 88.460 79.400 ;
        RECT 93.630 78.150 93.980 79.400 ;
        RECT 99.150 78.150 99.500 79.400 ;
        RECT 104.670 78.150 105.020 79.400 ;
        RECT 106.785 78.745 109.375 79.835 ;
        RECT 108.165 78.225 109.375 78.745 ;
        RECT 110.005 78.670 110.295 79.835 ;
        RECT 110.465 79.400 115.810 79.835 ;
        RECT 115.985 79.400 121.330 79.835 ;
        RECT 121.505 79.400 126.850 79.835 ;
        RECT 127.025 79.400 132.370 79.835 ;
        RECT 113.870 78.150 114.220 79.400 ;
        RECT 119.390 78.150 119.740 79.400 ;
        RECT 124.910 78.150 125.260 79.400 ;
        RECT 130.430 78.150 130.780 79.400 ;
        RECT 133.005 78.745 134.215 79.835 ;
        RECT 133.005 78.205 133.525 78.745 ;
        RECT 46.295 75.655 46.815 76.195 ;
        RECT 45.605 74.565 46.815 75.655 ;
        RECT 50.390 75.000 50.740 76.250 ;
        RECT 55.910 75.000 56.260 76.250 ;
        RECT 61.430 75.000 61.780 76.250 ;
        RECT 66.950 75.000 67.300 76.250 ;
        RECT 69.985 75.655 70.735 76.175 ;
        RECT 46.985 74.565 52.330 75.000 ;
        RECT 52.505 74.565 57.850 75.000 ;
        RECT 58.025 74.565 63.370 75.000 ;
        RECT 63.545 74.565 68.890 75.000 ;
        RECT 69.065 74.565 70.735 75.655 ;
        RECT 71.365 74.565 71.655 75.730 ;
        RECT 75.230 75.000 75.580 76.250 ;
        RECT 80.750 75.000 81.100 76.250 ;
        RECT 86.270 75.000 86.620 76.250 ;
        RECT 91.790 75.000 92.140 76.250 ;
        RECT 95.285 75.655 96.495 76.175 ;
        RECT 71.825 74.565 77.170 75.000 ;
        RECT 77.345 74.565 82.690 75.000 ;
        RECT 82.865 74.565 88.210 75.000 ;
        RECT 88.385 74.565 93.730 75.000 ;
        RECT 93.905 74.565 96.495 75.655 ;
        RECT 97.125 74.565 97.415 75.730 ;
        RECT 100.990 75.000 101.340 76.250 ;
        RECT 106.510 75.000 106.860 76.250 ;
        RECT 112.030 75.000 112.380 76.250 ;
        RECT 117.550 75.000 117.900 76.250 ;
        RECT 121.045 75.655 122.255 76.175 ;
        RECT 97.585 74.565 102.930 75.000 ;
        RECT 103.105 74.565 108.450 75.000 ;
        RECT 108.625 74.565 113.970 75.000 ;
        RECT 114.145 74.565 119.490 75.000 ;
        RECT 119.665 74.565 122.255 75.655 ;
        RECT 122.885 74.565 123.175 75.730 ;
        RECT 126.750 75.000 127.100 76.250 ;
        RECT 130.685 75.655 132.375 76.175 ;
        RECT 123.345 74.565 128.690 75.000 ;
        RECT 128.865 74.565 132.375 75.655 ;
        RECT 133.005 75.655 133.525 76.195 ;
        RECT 133.005 74.565 134.215 75.655 ;
        RECT 45.520 74.395 134.300 74.565 ;
        RECT 45.605 73.305 46.815 74.395 ;
        RECT 46.985 73.960 52.330 74.395 ;
        RECT 52.505 73.960 57.850 74.395 ;
        RECT 46.295 72.765 46.815 73.305 ;
        RECT 50.390 72.710 50.740 73.960 ;
        RECT 55.910 72.710 56.260 73.960 ;
        RECT 58.485 73.230 58.775 74.395 ;
        RECT 58.945 73.960 64.290 74.395 ;
        RECT 64.465 73.960 69.810 74.395 ;
        RECT 69.985 73.960 75.330 74.395 ;
        RECT 75.505 73.960 80.850 74.395 ;
        RECT 62.350 72.710 62.700 73.960 ;
        RECT 67.870 72.710 68.220 73.960 ;
        RECT 73.390 72.710 73.740 73.960 ;
        RECT 78.910 72.710 79.260 73.960 ;
        RECT 81.025 73.305 83.615 74.395 ;
        RECT 82.405 72.785 83.615 73.305 ;
        RECT 84.245 73.230 84.535 74.395 ;
        RECT 84.705 73.960 90.050 74.395 ;
        RECT 90.225 73.960 95.570 74.395 ;
        RECT 95.745 73.960 101.090 74.395 ;
        RECT 101.265 73.960 106.610 74.395 ;
        RECT 88.110 72.710 88.460 73.960 ;
        RECT 93.630 72.710 93.980 73.960 ;
        RECT 99.150 72.710 99.500 73.960 ;
        RECT 104.670 72.710 105.020 73.960 ;
        RECT 106.785 73.305 109.375 74.395 ;
        RECT 108.165 72.785 109.375 73.305 ;
        RECT 110.005 73.230 110.295 74.395 ;
        RECT 110.465 73.960 115.810 74.395 ;
        RECT 115.985 73.960 121.330 74.395 ;
        RECT 121.505 73.960 126.850 74.395 ;
        RECT 127.025 73.960 132.370 74.395 ;
        RECT 113.870 72.710 114.220 73.960 ;
        RECT 119.390 72.710 119.740 73.960 ;
        RECT 124.910 72.710 125.260 73.960 ;
        RECT 130.430 72.710 130.780 73.960 ;
        RECT 133.005 73.305 134.215 74.395 ;
        RECT 133.005 72.765 133.525 73.305 ;
        RECT 46.295 70.215 46.815 70.755 ;
        RECT 45.605 69.125 46.815 70.215 ;
        RECT 50.390 69.560 50.740 70.810 ;
        RECT 55.910 69.560 56.260 70.810 ;
        RECT 61.430 69.560 61.780 70.810 ;
        RECT 66.950 69.560 67.300 70.810 ;
        RECT 69.985 70.215 70.735 70.735 ;
        RECT 46.985 69.125 52.330 69.560 ;
        RECT 52.505 69.125 57.850 69.560 ;
        RECT 58.025 69.125 63.370 69.560 ;
        RECT 63.545 69.125 68.890 69.560 ;
        RECT 69.065 69.125 70.735 70.215 ;
        RECT 71.365 69.125 71.655 70.290 ;
        RECT 75.230 69.560 75.580 70.810 ;
        RECT 80.750 69.560 81.100 70.810 ;
        RECT 86.270 69.560 86.620 70.810 ;
        RECT 91.790 69.560 92.140 70.810 ;
        RECT 95.285 70.215 96.495 70.735 ;
        RECT 71.825 69.125 77.170 69.560 ;
        RECT 77.345 69.125 82.690 69.560 ;
        RECT 82.865 69.125 88.210 69.560 ;
        RECT 88.385 69.125 93.730 69.560 ;
        RECT 93.905 69.125 96.495 70.215 ;
        RECT 97.125 69.125 97.415 70.290 ;
        RECT 100.990 69.560 101.340 70.810 ;
        RECT 106.510 69.560 106.860 70.810 ;
        RECT 112.030 69.560 112.380 70.810 ;
        RECT 117.550 69.560 117.900 70.810 ;
        RECT 121.045 70.215 122.255 70.735 ;
        RECT 97.585 69.125 102.930 69.560 ;
        RECT 103.105 69.125 108.450 69.560 ;
        RECT 108.625 69.125 113.970 69.560 ;
        RECT 114.145 69.125 119.490 69.560 ;
        RECT 119.665 69.125 122.255 70.215 ;
        RECT 122.885 69.125 123.175 70.290 ;
        RECT 126.750 69.560 127.100 70.810 ;
        RECT 130.685 70.215 132.375 70.735 ;
        RECT 123.345 69.125 128.690 69.560 ;
        RECT 128.865 69.125 132.375 70.215 ;
        RECT 133.005 70.215 133.525 70.755 ;
        RECT 133.005 69.125 134.215 70.215 ;
        RECT 45.520 68.955 134.300 69.125 ;
        RECT 45.605 67.865 46.815 68.955 ;
        RECT 46.985 68.520 52.330 68.955 ;
        RECT 52.505 68.520 57.850 68.955 ;
        RECT 46.295 67.325 46.815 67.865 ;
        RECT 50.390 67.270 50.740 68.520 ;
        RECT 55.910 67.270 56.260 68.520 ;
        RECT 58.485 67.790 58.775 68.955 ;
        RECT 58.945 68.520 64.290 68.955 ;
        RECT 64.465 68.520 69.810 68.955 ;
        RECT 69.985 68.520 75.330 68.955 ;
        RECT 75.505 68.520 80.850 68.955 ;
        RECT 62.350 67.270 62.700 68.520 ;
        RECT 67.870 67.270 68.220 68.520 ;
        RECT 73.390 67.270 73.740 68.520 ;
        RECT 78.910 67.270 79.260 68.520 ;
        RECT 81.025 67.865 83.615 68.955 ;
        RECT 82.405 67.345 83.615 67.865 ;
        RECT 84.245 67.790 84.535 68.955 ;
        RECT 84.705 68.520 90.050 68.955 ;
        RECT 90.225 68.520 95.570 68.955 ;
        RECT 95.745 68.520 101.090 68.955 ;
        RECT 101.265 68.520 106.610 68.955 ;
        RECT 88.110 67.270 88.460 68.520 ;
        RECT 93.630 67.270 93.980 68.520 ;
        RECT 99.150 67.270 99.500 68.520 ;
        RECT 104.670 67.270 105.020 68.520 ;
        RECT 106.785 67.865 109.375 68.955 ;
        RECT 108.165 67.345 109.375 67.865 ;
        RECT 110.005 67.790 110.295 68.955 ;
        RECT 110.465 68.520 115.810 68.955 ;
        RECT 115.985 68.520 121.330 68.955 ;
        RECT 121.505 68.520 126.850 68.955 ;
        RECT 127.025 68.520 132.370 68.955 ;
        RECT 113.870 67.270 114.220 68.520 ;
        RECT 119.390 67.270 119.740 68.520 ;
        RECT 124.910 67.270 125.260 68.520 ;
        RECT 130.430 67.270 130.780 68.520 ;
        RECT 133.005 67.865 134.215 68.955 ;
        RECT 133.005 67.325 133.525 67.865 ;
        RECT 46.295 64.775 46.815 65.315 ;
        RECT 45.605 63.685 46.815 64.775 ;
        RECT 50.390 64.120 50.740 65.370 ;
        RECT 55.910 64.120 56.260 65.370 ;
        RECT 61.430 64.120 61.780 65.370 ;
        RECT 66.950 64.120 67.300 65.370 ;
        RECT 69.985 64.775 70.735 65.295 ;
        RECT 46.985 63.685 52.330 64.120 ;
        RECT 52.505 63.685 57.850 64.120 ;
        RECT 58.025 63.685 63.370 64.120 ;
        RECT 63.545 63.685 68.890 64.120 ;
        RECT 69.065 63.685 70.735 64.775 ;
        RECT 71.365 63.685 71.655 64.850 ;
        RECT 75.230 64.120 75.580 65.370 ;
        RECT 80.750 64.120 81.100 65.370 ;
        RECT 86.270 64.120 86.620 65.370 ;
        RECT 91.790 64.120 92.140 65.370 ;
        RECT 95.285 64.775 96.495 65.295 ;
        RECT 71.825 63.685 77.170 64.120 ;
        RECT 77.345 63.685 82.690 64.120 ;
        RECT 82.865 63.685 88.210 64.120 ;
        RECT 88.385 63.685 93.730 64.120 ;
        RECT 93.905 63.685 96.495 64.775 ;
        RECT 97.125 63.685 97.415 64.850 ;
        RECT 100.990 64.120 101.340 65.370 ;
        RECT 106.510 64.120 106.860 65.370 ;
        RECT 112.030 64.120 112.380 65.370 ;
        RECT 117.550 64.120 117.900 65.370 ;
        RECT 121.045 64.775 122.255 65.295 ;
        RECT 97.585 63.685 102.930 64.120 ;
        RECT 103.105 63.685 108.450 64.120 ;
        RECT 108.625 63.685 113.970 64.120 ;
        RECT 114.145 63.685 119.490 64.120 ;
        RECT 119.665 63.685 122.255 64.775 ;
        RECT 122.885 63.685 123.175 64.850 ;
        RECT 126.750 64.120 127.100 65.370 ;
        RECT 130.685 64.775 132.375 65.295 ;
        RECT 123.345 63.685 128.690 64.120 ;
        RECT 128.865 63.685 132.375 64.775 ;
        RECT 133.005 64.775 133.525 65.315 ;
        RECT 133.005 63.685 134.215 64.775 ;
        RECT 45.520 63.515 134.300 63.685 ;
        RECT 45.605 62.425 46.815 63.515 ;
        RECT 46.985 63.080 52.330 63.515 ;
        RECT 52.505 63.080 57.850 63.515 ;
        RECT 46.295 61.885 46.815 62.425 ;
        RECT 50.390 61.830 50.740 63.080 ;
        RECT 55.910 61.830 56.260 63.080 ;
        RECT 58.485 62.350 58.775 63.515 ;
        RECT 58.945 63.080 64.290 63.515 ;
        RECT 64.465 63.080 69.810 63.515 ;
        RECT 62.350 61.830 62.700 63.080 ;
        RECT 67.870 61.830 68.220 63.080 ;
        RECT 69.985 62.425 71.195 63.515 ;
        RECT 70.675 61.885 71.195 62.425 ;
        RECT 71.365 62.350 71.655 63.515 ;
        RECT 71.825 63.080 77.170 63.515 ;
        RECT 77.345 63.080 82.690 63.515 ;
        RECT 75.230 61.830 75.580 63.080 ;
        RECT 80.750 61.830 81.100 63.080 ;
        RECT 82.865 62.425 84.075 63.515 ;
        RECT 83.555 61.885 84.075 62.425 ;
        RECT 84.245 62.350 84.535 63.515 ;
        RECT 84.705 63.080 90.050 63.515 ;
        RECT 90.225 63.080 95.570 63.515 ;
        RECT 88.110 61.830 88.460 63.080 ;
        RECT 93.630 61.830 93.980 63.080 ;
        RECT 95.745 62.425 96.955 63.515 ;
        RECT 96.435 61.885 96.955 62.425 ;
        RECT 97.125 62.350 97.415 63.515 ;
        RECT 97.585 63.080 102.930 63.515 ;
        RECT 103.105 63.080 108.450 63.515 ;
        RECT 100.990 61.830 101.340 63.080 ;
        RECT 106.510 61.830 106.860 63.080 ;
        RECT 108.625 62.425 109.835 63.515 ;
        RECT 109.315 61.885 109.835 62.425 ;
        RECT 110.005 62.350 110.295 63.515 ;
        RECT 110.465 63.080 115.810 63.515 ;
        RECT 115.985 63.080 121.330 63.515 ;
        RECT 113.870 61.830 114.220 63.080 ;
        RECT 119.390 61.830 119.740 63.080 ;
        RECT 121.505 62.425 122.715 63.515 ;
        RECT 122.195 61.885 122.715 62.425 ;
        RECT 122.885 62.350 123.175 63.515 ;
        RECT 123.345 63.080 128.690 63.515 ;
        RECT 126.750 61.830 127.100 63.080 ;
        RECT 128.865 62.425 132.375 63.515 ;
        RECT 130.685 61.905 132.375 62.425 ;
        RECT 133.005 62.425 134.215 63.515 ;
        RECT 133.005 61.885 133.525 62.425 ;
      LAYER mcon ;
        RECT 45.665 134.235 45.835 134.405 ;
        RECT 46.125 134.235 46.295 134.405 ;
        RECT 46.585 134.235 46.755 134.405 ;
        RECT 47.045 134.235 47.215 134.405 ;
        RECT 47.505 134.235 47.675 134.405 ;
        RECT 47.965 134.235 48.135 134.405 ;
        RECT 48.425 134.235 48.595 134.405 ;
        RECT 48.885 134.235 49.055 134.405 ;
        RECT 49.345 134.235 49.515 134.405 ;
        RECT 49.805 134.235 49.975 134.405 ;
        RECT 50.265 134.235 50.435 134.405 ;
        RECT 50.725 134.235 50.895 134.405 ;
        RECT 51.185 134.235 51.355 134.405 ;
        RECT 51.645 134.235 51.815 134.405 ;
        RECT 52.105 134.235 52.275 134.405 ;
        RECT 52.565 134.235 52.735 134.405 ;
        RECT 53.025 134.235 53.195 134.405 ;
        RECT 53.485 134.235 53.655 134.405 ;
        RECT 53.945 134.235 54.115 134.405 ;
        RECT 54.405 134.235 54.575 134.405 ;
        RECT 54.865 134.235 55.035 134.405 ;
        RECT 55.325 134.235 55.495 134.405 ;
        RECT 55.785 134.235 55.955 134.405 ;
        RECT 56.245 134.235 56.415 134.405 ;
        RECT 56.705 134.235 56.875 134.405 ;
        RECT 57.165 134.235 57.335 134.405 ;
        RECT 57.625 134.235 57.795 134.405 ;
        RECT 58.085 134.235 58.255 134.405 ;
        RECT 58.545 134.235 58.715 134.405 ;
        RECT 59.005 134.235 59.175 134.405 ;
        RECT 59.465 134.235 59.635 134.405 ;
        RECT 59.925 134.235 60.095 134.405 ;
        RECT 60.385 134.235 60.555 134.405 ;
        RECT 60.845 134.235 61.015 134.405 ;
        RECT 61.305 134.235 61.475 134.405 ;
        RECT 61.765 134.235 61.935 134.405 ;
        RECT 62.225 134.235 62.395 134.405 ;
        RECT 62.685 134.235 62.855 134.405 ;
        RECT 63.145 134.235 63.315 134.405 ;
        RECT 63.605 134.235 63.775 134.405 ;
        RECT 64.065 134.235 64.235 134.405 ;
        RECT 64.525 134.235 64.695 134.405 ;
        RECT 64.985 134.235 65.155 134.405 ;
        RECT 65.445 134.235 65.615 134.405 ;
        RECT 65.905 134.235 66.075 134.405 ;
        RECT 66.365 134.235 66.535 134.405 ;
        RECT 66.825 134.235 66.995 134.405 ;
        RECT 67.285 134.235 67.455 134.405 ;
        RECT 67.745 134.235 67.915 134.405 ;
        RECT 68.205 134.235 68.375 134.405 ;
        RECT 68.665 134.235 68.835 134.405 ;
        RECT 69.125 134.235 69.295 134.405 ;
        RECT 69.585 134.235 69.755 134.405 ;
        RECT 70.045 134.235 70.215 134.405 ;
        RECT 70.505 134.235 70.675 134.405 ;
        RECT 70.965 134.235 71.135 134.405 ;
        RECT 71.425 134.235 71.595 134.405 ;
        RECT 71.885 134.235 72.055 134.405 ;
        RECT 72.345 134.235 72.515 134.405 ;
        RECT 72.805 134.235 72.975 134.405 ;
        RECT 73.265 134.235 73.435 134.405 ;
        RECT 73.725 134.235 73.895 134.405 ;
        RECT 74.185 134.235 74.355 134.405 ;
        RECT 74.645 134.235 74.815 134.405 ;
        RECT 75.105 134.235 75.275 134.405 ;
        RECT 75.565 134.235 75.735 134.405 ;
        RECT 76.025 134.235 76.195 134.405 ;
        RECT 76.485 134.235 76.655 134.405 ;
        RECT 76.945 134.235 77.115 134.405 ;
        RECT 77.405 134.235 77.575 134.405 ;
        RECT 77.865 134.235 78.035 134.405 ;
        RECT 78.325 134.235 78.495 134.405 ;
        RECT 78.785 134.235 78.955 134.405 ;
        RECT 79.245 134.235 79.415 134.405 ;
        RECT 79.705 134.235 79.875 134.405 ;
        RECT 80.165 134.235 80.335 134.405 ;
        RECT 80.625 134.235 80.795 134.405 ;
        RECT 81.085 134.235 81.255 134.405 ;
        RECT 81.545 134.235 81.715 134.405 ;
        RECT 82.005 134.235 82.175 134.405 ;
        RECT 82.465 134.235 82.635 134.405 ;
        RECT 82.925 134.235 83.095 134.405 ;
        RECT 83.385 134.235 83.555 134.405 ;
        RECT 83.845 134.235 84.015 134.405 ;
        RECT 84.305 134.235 84.475 134.405 ;
        RECT 84.765 134.235 84.935 134.405 ;
        RECT 85.225 134.235 85.395 134.405 ;
        RECT 85.685 134.235 85.855 134.405 ;
        RECT 86.145 134.235 86.315 134.405 ;
        RECT 86.605 134.235 86.775 134.405 ;
        RECT 87.065 134.235 87.235 134.405 ;
        RECT 87.525 134.235 87.695 134.405 ;
        RECT 87.985 134.235 88.155 134.405 ;
        RECT 88.445 134.235 88.615 134.405 ;
        RECT 88.905 134.235 89.075 134.405 ;
        RECT 89.365 134.235 89.535 134.405 ;
        RECT 89.825 134.235 89.995 134.405 ;
        RECT 90.285 134.235 90.455 134.405 ;
        RECT 90.745 134.235 90.915 134.405 ;
        RECT 91.205 134.235 91.375 134.405 ;
        RECT 91.665 134.235 91.835 134.405 ;
        RECT 92.125 134.235 92.295 134.405 ;
        RECT 92.585 134.235 92.755 134.405 ;
        RECT 93.045 134.235 93.215 134.405 ;
        RECT 93.505 134.235 93.675 134.405 ;
        RECT 93.965 134.235 94.135 134.405 ;
        RECT 94.425 134.235 94.595 134.405 ;
        RECT 94.885 134.235 95.055 134.405 ;
        RECT 95.345 134.235 95.515 134.405 ;
        RECT 95.805 134.235 95.975 134.405 ;
        RECT 96.265 134.235 96.435 134.405 ;
        RECT 96.725 134.235 96.895 134.405 ;
        RECT 97.185 134.235 97.355 134.405 ;
        RECT 97.645 134.235 97.815 134.405 ;
        RECT 98.105 134.235 98.275 134.405 ;
        RECT 98.565 134.235 98.735 134.405 ;
        RECT 99.025 134.235 99.195 134.405 ;
        RECT 99.485 134.235 99.655 134.405 ;
        RECT 99.945 134.235 100.115 134.405 ;
        RECT 100.405 134.235 100.575 134.405 ;
        RECT 100.865 134.235 101.035 134.405 ;
        RECT 101.325 134.235 101.495 134.405 ;
        RECT 101.785 134.235 101.955 134.405 ;
        RECT 102.245 134.235 102.415 134.405 ;
        RECT 102.705 134.235 102.875 134.405 ;
        RECT 103.165 134.235 103.335 134.405 ;
        RECT 103.625 134.235 103.795 134.405 ;
        RECT 104.085 134.235 104.255 134.405 ;
        RECT 104.545 134.235 104.715 134.405 ;
        RECT 105.005 134.235 105.175 134.405 ;
        RECT 105.465 134.235 105.635 134.405 ;
        RECT 105.925 134.235 106.095 134.405 ;
        RECT 106.385 134.235 106.555 134.405 ;
        RECT 106.845 134.235 107.015 134.405 ;
        RECT 107.305 134.235 107.475 134.405 ;
        RECT 107.765 134.235 107.935 134.405 ;
        RECT 108.225 134.235 108.395 134.405 ;
        RECT 108.685 134.235 108.855 134.405 ;
        RECT 109.145 134.235 109.315 134.405 ;
        RECT 109.605 134.235 109.775 134.405 ;
        RECT 110.065 134.235 110.235 134.405 ;
        RECT 110.525 134.235 110.695 134.405 ;
        RECT 110.985 134.235 111.155 134.405 ;
        RECT 111.445 134.235 111.615 134.405 ;
        RECT 111.905 134.235 112.075 134.405 ;
        RECT 112.365 134.235 112.535 134.405 ;
        RECT 112.825 134.235 112.995 134.405 ;
        RECT 113.285 134.235 113.455 134.405 ;
        RECT 113.745 134.235 113.915 134.405 ;
        RECT 114.205 134.235 114.375 134.405 ;
        RECT 114.665 134.235 114.835 134.405 ;
        RECT 115.125 134.235 115.295 134.405 ;
        RECT 115.585 134.235 115.755 134.405 ;
        RECT 116.045 134.235 116.215 134.405 ;
        RECT 116.505 134.235 116.675 134.405 ;
        RECT 116.965 134.235 117.135 134.405 ;
        RECT 117.425 134.235 117.595 134.405 ;
        RECT 117.885 134.235 118.055 134.405 ;
        RECT 118.345 134.235 118.515 134.405 ;
        RECT 118.805 134.235 118.975 134.405 ;
        RECT 119.265 134.235 119.435 134.405 ;
        RECT 119.725 134.235 119.895 134.405 ;
        RECT 120.185 134.235 120.355 134.405 ;
        RECT 120.645 134.235 120.815 134.405 ;
        RECT 121.105 134.235 121.275 134.405 ;
        RECT 121.565 134.235 121.735 134.405 ;
        RECT 122.025 134.235 122.195 134.405 ;
        RECT 122.485 134.235 122.655 134.405 ;
        RECT 122.945 134.235 123.115 134.405 ;
        RECT 123.405 134.235 123.575 134.405 ;
        RECT 123.865 134.235 124.035 134.405 ;
        RECT 124.325 134.235 124.495 134.405 ;
        RECT 124.785 134.235 124.955 134.405 ;
        RECT 125.245 134.235 125.415 134.405 ;
        RECT 125.705 134.235 125.875 134.405 ;
        RECT 126.165 134.235 126.335 134.405 ;
        RECT 126.625 134.235 126.795 134.405 ;
        RECT 127.085 134.235 127.255 134.405 ;
        RECT 127.545 134.235 127.715 134.405 ;
        RECT 128.005 134.235 128.175 134.405 ;
        RECT 128.465 134.235 128.635 134.405 ;
        RECT 128.925 134.235 129.095 134.405 ;
        RECT 129.385 134.235 129.555 134.405 ;
        RECT 129.845 134.235 130.015 134.405 ;
        RECT 130.305 134.235 130.475 134.405 ;
        RECT 130.765 134.235 130.935 134.405 ;
        RECT 131.225 134.235 131.395 134.405 ;
        RECT 131.685 134.235 131.855 134.405 ;
        RECT 132.145 134.235 132.315 134.405 ;
        RECT 132.605 134.235 132.775 134.405 ;
        RECT 133.065 134.235 133.235 134.405 ;
        RECT 133.525 134.235 133.695 134.405 ;
        RECT 133.985 134.235 134.155 134.405 ;
        RECT 45.665 128.795 45.835 128.965 ;
        RECT 46.125 128.795 46.295 128.965 ;
        RECT 46.585 128.795 46.755 128.965 ;
        RECT 47.045 128.795 47.215 128.965 ;
        RECT 47.505 128.795 47.675 128.965 ;
        RECT 47.965 128.795 48.135 128.965 ;
        RECT 48.425 128.795 48.595 128.965 ;
        RECT 48.885 128.795 49.055 128.965 ;
        RECT 49.345 128.795 49.515 128.965 ;
        RECT 49.805 128.795 49.975 128.965 ;
        RECT 50.265 128.795 50.435 128.965 ;
        RECT 50.725 128.795 50.895 128.965 ;
        RECT 51.185 128.795 51.355 128.965 ;
        RECT 51.645 128.795 51.815 128.965 ;
        RECT 52.105 128.795 52.275 128.965 ;
        RECT 52.565 128.795 52.735 128.965 ;
        RECT 53.025 128.795 53.195 128.965 ;
        RECT 53.485 128.795 53.655 128.965 ;
        RECT 53.945 128.795 54.115 128.965 ;
        RECT 54.405 128.795 54.575 128.965 ;
        RECT 54.865 128.795 55.035 128.965 ;
        RECT 55.325 128.795 55.495 128.965 ;
        RECT 55.785 128.795 55.955 128.965 ;
        RECT 56.245 128.795 56.415 128.965 ;
        RECT 56.705 128.795 56.875 128.965 ;
        RECT 57.165 128.795 57.335 128.965 ;
        RECT 57.625 128.795 57.795 128.965 ;
        RECT 58.085 128.795 58.255 128.965 ;
        RECT 58.545 128.795 58.715 128.965 ;
        RECT 59.005 128.795 59.175 128.965 ;
        RECT 59.465 128.795 59.635 128.965 ;
        RECT 59.925 128.795 60.095 128.965 ;
        RECT 60.385 128.795 60.555 128.965 ;
        RECT 60.845 128.795 61.015 128.965 ;
        RECT 61.305 128.795 61.475 128.965 ;
        RECT 61.765 128.795 61.935 128.965 ;
        RECT 62.225 128.795 62.395 128.965 ;
        RECT 62.685 128.795 62.855 128.965 ;
        RECT 63.145 128.795 63.315 128.965 ;
        RECT 63.605 128.795 63.775 128.965 ;
        RECT 64.065 128.795 64.235 128.965 ;
        RECT 64.525 128.795 64.695 128.965 ;
        RECT 64.985 128.795 65.155 128.965 ;
        RECT 65.445 128.795 65.615 128.965 ;
        RECT 65.905 128.795 66.075 128.965 ;
        RECT 66.365 128.795 66.535 128.965 ;
        RECT 66.825 128.795 66.995 128.965 ;
        RECT 67.285 128.795 67.455 128.965 ;
        RECT 67.745 128.795 67.915 128.965 ;
        RECT 68.205 128.795 68.375 128.965 ;
        RECT 68.665 128.795 68.835 128.965 ;
        RECT 69.125 128.795 69.295 128.965 ;
        RECT 69.585 128.795 69.755 128.965 ;
        RECT 70.045 128.795 70.215 128.965 ;
        RECT 70.505 128.795 70.675 128.965 ;
        RECT 70.965 128.795 71.135 128.965 ;
        RECT 71.425 128.795 71.595 128.965 ;
        RECT 71.885 128.795 72.055 128.965 ;
        RECT 72.345 128.795 72.515 128.965 ;
        RECT 72.805 128.795 72.975 128.965 ;
        RECT 73.265 128.795 73.435 128.965 ;
        RECT 73.725 128.795 73.895 128.965 ;
        RECT 74.185 128.795 74.355 128.965 ;
        RECT 74.645 128.795 74.815 128.965 ;
        RECT 75.105 128.795 75.275 128.965 ;
        RECT 75.565 128.795 75.735 128.965 ;
        RECT 76.025 128.795 76.195 128.965 ;
        RECT 76.485 128.795 76.655 128.965 ;
        RECT 76.945 128.795 77.115 128.965 ;
        RECT 77.405 128.795 77.575 128.965 ;
        RECT 77.865 128.795 78.035 128.965 ;
        RECT 78.325 128.795 78.495 128.965 ;
        RECT 78.785 128.795 78.955 128.965 ;
        RECT 79.245 128.795 79.415 128.965 ;
        RECT 79.705 128.795 79.875 128.965 ;
        RECT 80.165 128.795 80.335 128.965 ;
        RECT 80.625 128.795 80.795 128.965 ;
        RECT 81.085 128.795 81.255 128.965 ;
        RECT 81.545 128.795 81.715 128.965 ;
        RECT 82.005 128.795 82.175 128.965 ;
        RECT 82.465 128.795 82.635 128.965 ;
        RECT 82.925 128.795 83.095 128.965 ;
        RECT 83.385 128.795 83.555 128.965 ;
        RECT 83.845 128.795 84.015 128.965 ;
        RECT 84.305 128.795 84.475 128.965 ;
        RECT 84.765 128.795 84.935 128.965 ;
        RECT 85.225 128.795 85.395 128.965 ;
        RECT 85.685 128.795 85.855 128.965 ;
        RECT 86.145 128.795 86.315 128.965 ;
        RECT 86.605 128.795 86.775 128.965 ;
        RECT 87.065 128.795 87.235 128.965 ;
        RECT 87.525 128.795 87.695 128.965 ;
        RECT 87.985 128.795 88.155 128.965 ;
        RECT 88.445 128.795 88.615 128.965 ;
        RECT 88.905 128.795 89.075 128.965 ;
        RECT 89.365 128.795 89.535 128.965 ;
        RECT 89.825 128.795 89.995 128.965 ;
        RECT 90.285 128.795 90.455 128.965 ;
        RECT 90.745 128.795 90.915 128.965 ;
        RECT 91.205 128.795 91.375 128.965 ;
        RECT 91.665 128.795 91.835 128.965 ;
        RECT 92.125 128.795 92.295 128.965 ;
        RECT 92.585 128.795 92.755 128.965 ;
        RECT 93.045 128.795 93.215 128.965 ;
        RECT 93.505 128.795 93.675 128.965 ;
        RECT 93.965 128.795 94.135 128.965 ;
        RECT 94.425 128.795 94.595 128.965 ;
        RECT 94.885 128.795 95.055 128.965 ;
        RECT 95.345 128.795 95.515 128.965 ;
        RECT 95.805 128.795 95.975 128.965 ;
        RECT 96.265 128.795 96.435 128.965 ;
        RECT 96.725 128.795 96.895 128.965 ;
        RECT 97.185 128.795 97.355 128.965 ;
        RECT 97.645 128.795 97.815 128.965 ;
        RECT 98.105 128.795 98.275 128.965 ;
        RECT 98.565 128.795 98.735 128.965 ;
        RECT 99.025 128.795 99.195 128.965 ;
        RECT 99.485 128.795 99.655 128.965 ;
        RECT 99.945 128.795 100.115 128.965 ;
        RECT 100.405 128.795 100.575 128.965 ;
        RECT 100.865 128.795 101.035 128.965 ;
        RECT 101.325 128.795 101.495 128.965 ;
        RECT 101.785 128.795 101.955 128.965 ;
        RECT 102.245 128.795 102.415 128.965 ;
        RECT 102.705 128.795 102.875 128.965 ;
        RECT 103.165 128.795 103.335 128.965 ;
        RECT 103.625 128.795 103.795 128.965 ;
        RECT 104.085 128.795 104.255 128.965 ;
        RECT 104.545 128.795 104.715 128.965 ;
        RECT 105.005 128.795 105.175 128.965 ;
        RECT 105.465 128.795 105.635 128.965 ;
        RECT 105.925 128.795 106.095 128.965 ;
        RECT 106.385 128.795 106.555 128.965 ;
        RECT 106.845 128.795 107.015 128.965 ;
        RECT 107.305 128.795 107.475 128.965 ;
        RECT 107.765 128.795 107.935 128.965 ;
        RECT 108.225 128.795 108.395 128.965 ;
        RECT 108.685 128.795 108.855 128.965 ;
        RECT 109.145 128.795 109.315 128.965 ;
        RECT 109.605 128.795 109.775 128.965 ;
        RECT 110.065 128.795 110.235 128.965 ;
        RECT 110.525 128.795 110.695 128.965 ;
        RECT 110.985 128.795 111.155 128.965 ;
        RECT 111.445 128.795 111.615 128.965 ;
        RECT 111.905 128.795 112.075 128.965 ;
        RECT 112.365 128.795 112.535 128.965 ;
        RECT 112.825 128.795 112.995 128.965 ;
        RECT 113.285 128.795 113.455 128.965 ;
        RECT 113.745 128.795 113.915 128.965 ;
        RECT 114.205 128.795 114.375 128.965 ;
        RECT 114.665 128.795 114.835 128.965 ;
        RECT 115.125 128.795 115.295 128.965 ;
        RECT 115.585 128.795 115.755 128.965 ;
        RECT 116.045 128.795 116.215 128.965 ;
        RECT 116.505 128.795 116.675 128.965 ;
        RECT 116.965 128.795 117.135 128.965 ;
        RECT 117.425 128.795 117.595 128.965 ;
        RECT 117.885 128.795 118.055 128.965 ;
        RECT 118.345 128.795 118.515 128.965 ;
        RECT 118.805 128.795 118.975 128.965 ;
        RECT 119.265 128.795 119.435 128.965 ;
        RECT 119.725 128.795 119.895 128.965 ;
        RECT 120.185 128.795 120.355 128.965 ;
        RECT 120.645 128.795 120.815 128.965 ;
        RECT 121.105 128.795 121.275 128.965 ;
        RECT 121.565 128.795 121.735 128.965 ;
        RECT 122.025 128.795 122.195 128.965 ;
        RECT 122.485 128.795 122.655 128.965 ;
        RECT 122.945 128.795 123.115 128.965 ;
        RECT 123.405 128.795 123.575 128.965 ;
        RECT 123.865 128.795 124.035 128.965 ;
        RECT 124.325 128.795 124.495 128.965 ;
        RECT 124.785 128.795 124.955 128.965 ;
        RECT 125.245 128.795 125.415 128.965 ;
        RECT 125.705 128.795 125.875 128.965 ;
        RECT 126.165 128.795 126.335 128.965 ;
        RECT 126.625 128.795 126.795 128.965 ;
        RECT 127.085 128.795 127.255 128.965 ;
        RECT 127.545 128.795 127.715 128.965 ;
        RECT 128.005 128.795 128.175 128.965 ;
        RECT 128.465 128.795 128.635 128.965 ;
        RECT 128.925 128.795 129.095 128.965 ;
        RECT 129.385 128.795 129.555 128.965 ;
        RECT 129.845 128.795 130.015 128.965 ;
        RECT 130.305 128.795 130.475 128.965 ;
        RECT 130.765 128.795 130.935 128.965 ;
        RECT 131.225 128.795 131.395 128.965 ;
        RECT 131.685 128.795 131.855 128.965 ;
        RECT 132.145 128.795 132.315 128.965 ;
        RECT 132.605 128.795 132.775 128.965 ;
        RECT 133.065 128.795 133.235 128.965 ;
        RECT 133.525 128.795 133.695 128.965 ;
        RECT 133.985 128.795 134.155 128.965 ;
        RECT 45.665 123.355 45.835 123.525 ;
        RECT 46.125 123.355 46.295 123.525 ;
        RECT 46.585 123.355 46.755 123.525 ;
        RECT 47.045 123.355 47.215 123.525 ;
        RECT 47.505 123.355 47.675 123.525 ;
        RECT 47.965 123.355 48.135 123.525 ;
        RECT 48.425 123.355 48.595 123.525 ;
        RECT 48.885 123.355 49.055 123.525 ;
        RECT 49.345 123.355 49.515 123.525 ;
        RECT 49.805 123.355 49.975 123.525 ;
        RECT 50.265 123.355 50.435 123.525 ;
        RECT 50.725 123.355 50.895 123.525 ;
        RECT 51.185 123.355 51.355 123.525 ;
        RECT 51.645 123.355 51.815 123.525 ;
        RECT 52.105 123.355 52.275 123.525 ;
        RECT 52.565 123.355 52.735 123.525 ;
        RECT 53.025 123.355 53.195 123.525 ;
        RECT 53.485 123.355 53.655 123.525 ;
        RECT 53.945 123.355 54.115 123.525 ;
        RECT 54.405 123.355 54.575 123.525 ;
        RECT 54.865 123.355 55.035 123.525 ;
        RECT 55.325 123.355 55.495 123.525 ;
        RECT 55.785 123.355 55.955 123.525 ;
        RECT 56.245 123.355 56.415 123.525 ;
        RECT 56.705 123.355 56.875 123.525 ;
        RECT 57.165 123.355 57.335 123.525 ;
        RECT 57.625 123.355 57.795 123.525 ;
        RECT 58.085 123.355 58.255 123.525 ;
        RECT 58.545 123.355 58.715 123.525 ;
        RECT 59.005 123.355 59.175 123.525 ;
        RECT 59.465 123.355 59.635 123.525 ;
        RECT 59.925 123.355 60.095 123.525 ;
        RECT 60.385 123.355 60.555 123.525 ;
        RECT 60.845 123.355 61.015 123.525 ;
        RECT 61.305 123.355 61.475 123.525 ;
        RECT 61.765 123.355 61.935 123.525 ;
        RECT 62.225 123.355 62.395 123.525 ;
        RECT 62.685 123.355 62.855 123.525 ;
        RECT 63.145 123.355 63.315 123.525 ;
        RECT 63.605 123.355 63.775 123.525 ;
        RECT 64.065 123.355 64.235 123.525 ;
        RECT 64.525 123.355 64.695 123.525 ;
        RECT 64.985 123.355 65.155 123.525 ;
        RECT 65.445 123.355 65.615 123.525 ;
        RECT 65.905 123.355 66.075 123.525 ;
        RECT 66.365 123.355 66.535 123.525 ;
        RECT 66.825 123.355 66.995 123.525 ;
        RECT 67.285 123.355 67.455 123.525 ;
        RECT 67.745 123.355 67.915 123.525 ;
        RECT 68.205 123.355 68.375 123.525 ;
        RECT 68.665 123.355 68.835 123.525 ;
        RECT 69.125 123.355 69.295 123.525 ;
        RECT 69.585 123.355 69.755 123.525 ;
        RECT 70.045 123.355 70.215 123.525 ;
        RECT 70.505 123.355 70.675 123.525 ;
        RECT 70.965 123.355 71.135 123.525 ;
        RECT 71.425 123.355 71.595 123.525 ;
        RECT 71.885 123.355 72.055 123.525 ;
        RECT 72.345 123.355 72.515 123.525 ;
        RECT 72.805 123.355 72.975 123.525 ;
        RECT 73.265 123.355 73.435 123.525 ;
        RECT 73.725 123.355 73.895 123.525 ;
        RECT 74.185 123.355 74.355 123.525 ;
        RECT 74.645 123.355 74.815 123.525 ;
        RECT 75.105 123.355 75.275 123.525 ;
        RECT 75.565 123.355 75.735 123.525 ;
        RECT 76.025 123.355 76.195 123.525 ;
        RECT 76.485 123.355 76.655 123.525 ;
        RECT 76.945 123.355 77.115 123.525 ;
        RECT 77.405 123.355 77.575 123.525 ;
        RECT 77.865 123.355 78.035 123.525 ;
        RECT 78.325 123.355 78.495 123.525 ;
        RECT 78.785 123.355 78.955 123.525 ;
        RECT 79.245 123.355 79.415 123.525 ;
        RECT 79.705 123.355 79.875 123.525 ;
        RECT 80.165 123.355 80.335 123.525 ;
        RECT 80.625 123.355 80.795 123.525 ;
        RECT 81.085 123.355 81.255 123.525 ;
        RECT 81.545 123.355 81.715 123.525 ;
        RECT 82.005 123.355 82.175 123.525 ;
        RECT 82.465 123.355 82.635 123.525 ;
        RECT 82.925 123.355 83.095 123.525 ;
        RECT 83.385 123.355 83.555 123.525 ;
        RECT 83.845 123.355 84.015 123.525 ;
        RECT 84.305 123.355 84.475 123.525 ;
        RECT 84.765 123.355 84.935 123.525 ;
        RECT 85.225 123.355 85.395 123.525 ;
        RECT 85.685 123.355 85.855 123.525 ;
        RECT 86.145 123.355 86.315 123.525 ;
        RECT 86.605 123.355 86.775 123.525 ;
        RECT 87.065 123.355 87.235 123.525 ;
        RECT 87.525 123.355 87.695 123.525 ;
        RECT 87.985 123.355 88.155 123.525 ;
        RECT 88.445 123.355 88.615 123.525 ;
        RECT 88.905 123.355 89.075 123.525 ;
        RECT 89.365 123.355 89.535 123.525 ;
        RECT 89.825 123.355 89.995 123.525 ;
        RECT 90.285 123.355 90.455 123.525 ;
        RECT 90.745 123.355 90.915 123.525 ;
        RECT 91.205 123.355 91.375 123.525 ;
        RECT 91.665 123.355 91.835 123.525 ;
        RECT 92.125 123.355 92.295 123.525 ;
        RECT 92.585 123.355 92.755 123.525 ;
        RECT 93.045 123.355 93.215 123.525 ;
        RECT 93.505 123.355 93.675 123.525 ;
        RECT 93.965 123.355 94.135 123.525 ;
        RECT 94.425 123.355 94.595 123.525 ;
        RECT 94.885 123.355 95.055 123.525 ;
        RECT 95.345 123.355 95.515 123.525 ;
        RECT 95.805 123.355 95.975 123.525 ;
        RECT 96.265 123.355 96.435 123.525 ;
        RECT 96.725 123.355 96.895 123.525 ;
        RECT 97.185 123.355 97.355 123.525 ;
        RECT 97.645 123.355 97.815 123.525 ;
        RECT 98.105 123.355 98.275 123.525 ;
        RECT 98.565 123.355 98.735 123.525 ;
        RECT 99.025 123.355 99.195 123.525 ;
        RECT 99.485 123.355 99.655 123.525 ;
        RECT 99.945 123.355 100.115 123.525 ;
        RECT 100.405 123.355 100.575 123.525 ;
        RECT 100.865 123.355 101.035 123.525 ;
        RECT 101.325 123.355 101.495 123.525 ;
        RECT 101.785 123.355 101.955 123.525 ;
        RECT 102.245 123.355 102.415 123.525 ;
        RECT 102.705 123.355 102.875 123.525 ;
        RECT 103.165 123.355 103.335 123.525 ;
        RECT 103.625 123.355 103.795 123.525 ;
        RECT 104.085 123.355 104.255 123.525 ;
        RECT 104.545 123.355 104.715 123.525 ;
        RECT 105.005 123.355 105.175 123.525 ;
        RECT 105.465 123.355 105.635 123.525 ;
        RECT 105.925 123.355 106.095 123.525 ;
        RECT 106.385 123.355 106.555 123.525 ;
        RECT 106.845 123.355 107.015 123.525 ;
        RECT 107.305 123.355 107.475 123.525 ;
        RECT 107.765 123.355 107.935 123.525 ;
        RECT 108.225 123.355 108.395 123.525 ;
        RECT 108.685 123.355 108.855 123.525 ;
        RECT 109.145 123.355 109.315 123.525 ;
        RECT 109.605 123.355 109.775 123.525 ;
        RECT 110.065 123.355 110.235 123.525 ;
        RECT 110.525 123.355 110.695 123.525 ;
        RECT 110.985 123.355 111.155 123.525 ;
        RECT 111.445 123.355 111.615 123.525 ;
        RECT 111.905 123.355 112.075 123.525 ;
        RECT 112.365 123.355 112.535 123.525 ;
        RECT 112.825 123.355 112.995 123.525 ;
        RECT 113.285 123.355 113.455 123.525 ;
        RECT 113.745 123.355 113.915 123.525 ;
        RECT 114.205 123.355 114.375 123.525 ;
        RECT 114.665 123.355 114.835 123.525 ;
        RECT 115.125 123.355 115.295 123.525 ;
        RECT 115.585 123.355 115.755 123.525 ;
        RECT 116.045 123.355 116.215 123.525 ;
        RECT 116.505 123.355 116.675 123.525 ;
        RECT 116.965 123.355 117.135 123.525 ;
        RECT 117.425 123.355 117.595 123.525 ;
        RECT 117.885 123.355 118.055 123.525 ;
        RECT 118.345 123.355 118.515 123.525 ;
        RECT 118.805 123.355 118.975 123.525 ;
        RECT 119.265 123.355 119.435 123.525 ;
        RECT 119.725 123.355 119.895 123.525 ;
        RECT 120.185 123.355 120.355 123.525 ;
        RECT 120.645 123.355 120.815 123.525 ;
        RECT 121.105 123.355 121.275 123.525 ;
        RECT 121.565 123.355 121.735 123.525 ;
        RECT 122.025 123.355 122.195 123.525 ;
        RECT 122.485 123.355 122.655 123.525 ;
        RECT 122.945 123.355 123.115 123.525 ;
        RECT 123.405 123.355 123.575 123.525 ;
        RECT 123.865 123.355 124.035 123.525 ;
        RECT 124.325 123.355 124.495 123.525 ;
        RECT 124.785 123.355 124.955 123.525 ;
        RECT 125.245 123.355 125.415 123.525 ;
        RECT 125.705 123.355 125.875 123.525 ;
        RECT 126.165 123.355 126.335 123.525 ;
        RECT 126.625 123.355 126.795 123.525 ;
        RECT 127.085 123.355 127.255 123.525 ;
        RECT 127.545 123.355 127.715 123.525 ;
        RECT 128.005 123.355 128.175 123.525 ;
        RECT 128.465 123.355 128.635 123.525 ;
        RECT 128.925 123.355 129.095 123.525 ;
        RECT 129.385 123.355 129.555 123.525 ;
        RECT 129.845 123.355 130.015 123.525 ;
        RECT 130.305 123.355 130.475 123.525 ;
        RECT 130.765 123.355 130.935 123.525 ;
        RECT 131.225 123.355 131.395 123.525 ;
        RECT 131.685 123.355 131.855 123.525 ;
        RECT 132.145 123.355 132.315 123.525 ;
        RECT 132.605 123.355 132.775 123.525 ;
        RECT 133.065 123.355 133.235 123.525 ;
        RECT 133.525 123.355 133.695 123.525 ;
        RECT 133.985 123.355 134.155 123.525 ;
        RECT 45.665 117.915 45.835 118.085 ;
        RECT 46.125 117.915 46.295 118.085 ;
        RECT 46.585 117.915 46.755 118.085 ;
        RECT 47.045 117.915 47.215 118.085 ;
        RECT 47.505 117.915 47.675 118.085 ;
        RECT 47.965 117.915 48.135 118.085 ;
        RECT 48.425 117.915 48.595 118.085 ;
        RECT 48.885 117.915 49.055 118.085 ;
        RECT 49.345 117.915 49.515 118.085 ;
        RECT 49.805 117.915 49.975 118.085 ;
        RECT 50.265 117.915 50.435 118.085 ;
        RECT 50.725 117.915 50.895 118.085 ;
        RECT 51.185 117.915 51.355 118.085 ;
        RECT 51.645 117.915 51.815 118.085 ;
        RECT 52.105 117.915 52.275 118.085 ;
        RECT 52.565 117.915 52.735 118.085 ;
        RECT 53.025 117.915 53.195 118.085 ;
        RECT 53.485 117.915 53.655 118.085 ;
        RECT 53.945 117.915 54.115 118.085 ;
        RECT 54.405 117.915 54.575 118.085 ;
        RECT 54.865 117.915 55.035 118.085 ;
        RECT 55.325 117.915 55.495 118.085 ;
        RECT 55.785 117.915 55.955 118.085 ;
        RECT 56.245 117.915 56.415 118.085 ;
        RECT 56.705 117.915 56.875 118.085 ;
        RECT 57.165 117.915 57.335 118.085 ;
        RECT 57.625 117.915 57.795 118.085 ;
        RECT 58.085 117.915 58.255 118.085 ;
        RECT 58.545 117.915 58.715 118.085 ;
        RECT 59.005 117.915 59.175 118.085 ;
        RECT 59.465 117.915 59.635 118.085 ;
        RECT 59.925 117.915 60.095 118.085 ;
        RECT 60.385 117.915 60.555 118.085 ;
        RECT 60.845 117.915 61.015 118.085 ;
        RECT 61.305 117.915 61.475 118.085 ;
        RECT 61.765 117.915 61.935 118.085 ;
        RECT 62.225 117.915 62.395 118.085 ;
        RECT 62.685 117.915 62.855 118.085 ;
        RECT 63.145 117.915 63.315 118.085 ;
        RECT 63.605 117.915 63.775 118.085 ;
        RECT 64.065 117.915 64.235 118.085 ;
        RECT 64.525 117.915 64.695 118.085 ;
        RECT 64.985 117.915 65.155 118.085 ;
        RECT 65.445 117.915 65.615 118.085 ;
        RECT 65.905 117.915 66.075 118.085 ;
        RECT 66.365 117.915 66.535 118.085 ;
        RECT 66.825 117.915 66.995 118.085 ;
        RECT 67.285 117.915 67.455 118.085 ;
        RECT 67.745 117.915 67.915 118.085 ;
        RECT 68.205 117.915 68.375 118.085 ;
        RECT 68.665 117.915 68.835 118.085 ;
        RECT 69.125 117.915 69.295 118.085 ;
        RECT 69.585 117.915 69.755 118.085 ;
        RECT 70.045 117.915 70.215 118.085 ;
        RECT 70.505 117.915 70.675 118.085 ;
        RECT 70.965 117.915 71.135 118.085 ;
        RECT 71.425 117.915 71.595 118.085 ;
        RECT 71.885 117.915 72.055 118.085 ;
        RECT 72.345 117.915 72.515 118.085 ;
        RECT 72.805 117.915 72.975 118.085 ;
        RECT 73.265 117.915 73.435 118.085 ;
        RECT 73.725 117.915 73.895 118.085 ;
        RECT 74.185 117.915 74.355 118.085 ;
        RECT 74.645 117.915 74.815 118.085 ;
        RECT 75.105 117.915 75.275 118.085 ;
        RECT 75.565 117.915 75.735 118.085 ;
        RECT 76.025 117.915 76.195 118.085 ;
        RECT 76.485 117.915 76.655 118.085 ;
        RECT 76.945 117.915 77.115 118.085 ;
        RECT 77.405 117.915 77.575 118.085 ;
        RECT 77.865 117.915 78.035 118.085 ;
        RECT 78.325 117.915 78.495 118.085 ;
        RECT 78.785 117.915 78.955 118.085 ;
        RECT 79.245 117.915 79.415 118.085 ;
        RECT 79.705 117.915 79.875 118.085 ;
        RECT 80.165 117.915 80.335 118.085 ;
        RECT 80.625 117.915 80.795 118.085 ;
        RECT 81.085 117.915 81.255 118.085 ;
        RECT 81.545 117.915 81.715 118.085 ;
        RECT 82.005 117.915 82.175 118.085 ;
        RECT 82.465 117.915 82.635 118.085 ;
        RECT 82.925 117.915 83.095 118.085 ;
        RECT 83.385 117.915 83.555 118.085 ;
        RECT 83.845 117.915 84.015 118.085 ;
        RECT 84.305 117.915 84.475 118.085 ;
        RECT 84.765 117.915 84.935 118.085 ;
        RECT 85.225 117.915 85.395 118.085 ;
        RECT 85.685 117.915 85.855 118.085 ;
        RECT 86.145 117.915 86.315 118.085 ;
        RECT 86.605 117.915 86.775 118.085 ;
        RECT 87.065 117.915 87.235 118.085 ;
        RECT 87.525 117.915 87.695 118.085 ;
        RECT 87.985 117.915 88.155 118.085 ;
        RECT 88.445 117.915 88.615 118.085 ;
        RECT 88.905 117.915 89.075 118.085 ;
        RECT 89.365 117.915 89.535 118.085 ;
        RECT 89.825 117.915 89.995 118.085 ;
        RECT 90.285 117.915 90.455 118.085 ;
        RECT 90.745 117.915 90.915 118.085 ;
        RECT 91.205 117.915 91.375 118.085 ;
        RECT 91.665 117.915 91.835 118.085 ;
        RECT 92.125 117.915 92.295 118.085 ;
        RECT 92.585 117.915 92.755 118.085 ;
        RECT 93.045 117.915 93.215 118.085 ;
        RECT 93.505 117.915 93.675 118.085 ;
        RECT 93.965 117.915 94.135 118.085 ;
        RECT 94.425 117.915 94.595 118.085 ;
        RECT 94.885 117.915 95.055 118.085 ;
        RECT 95.345 117.915 95.515 118.085 ;
        RECT 95.805 117.915 95.975 118.085 ;
        RECT 96.265 117.915 96.435 118.085 ;
        RECT 96.725 117.915 96.895 118.085 ;
        RECT 97.185 117.915 97.355 118.085 ;
        RECT 97.645 117.915 97.815 118.085 ;
        RECT 98.105 117.915 98.275 118.085 ;
        RECT 98.565 117.915 98.735 118.085 ;
        RECT 99.025 117.915 99.195 118.085 ;
        RECT 99.485 117.915 99.655 118.085 ;
        RECT 99.945 117.915 100.115 118.085 ;
        RECT 100.405 117.915 100.575 118.085 ;
        RECT 100.865 117.915 101.035 118.085 ;
        RECT 101.325 117.915 101.495 118.085 ;
        RECT 101.785 117.915 101.955 118.085 ;
        RECT 102.245 117.915 102.415 118.085 ;
        RECT 102.705 117.915 102.875 118.085 ;
        RECT 103.165 117.915 103.335 118.085 ;
        RECT 103.625 117.915 103.795 118.085 ;
        RECT 104.085 117.915 104.255 118.085 ;
        RECT 104.545 117.915 104.715 118.085 ;
        RECT 105.005 117.915 105.175 118.085 ;
        RECT 105.465 117.915 105.635 118.085 ;
        RECT 105.925 117.915 106.095 118.085 ;
        RECT 106.385 117.915 106.555 118.085 ;
        RECT 106.845 117.915 107.015 118.085 ;
        RECT 107.305 117.915 107.475 118.085 ;
        RECT 107.765 117.915 107.935 118.085 ;
        RECT 108.225 117.915 108.395 118.085 ;
        RECT 108.685 117.915 108.855 118.085 ;
        RECT 109.145 117.915 109.315 118.085 ;
        RECT 109.605 117.915 109.775 118.085 ;
        RECT 110.065 117.915 110.235 118.085 ;
        RECT 110.525 117.915 110.695 118.085 ;
        RECT 110.985 117.915 111.155 118.085 ;
        RECT 111.445 117.915 111.615 118.085 ;
        RECT 111.905 117.915 112.075 118.085 ;
        RECT 112.365 117.915 112.535 118.085 ;
        RECT 112.825 117.915 112.995 118.085 ;
        RECT 113.285 117.915 113.455 118.085 ;
        RECT 113.745 117.915 113.915 118.085 ;
        RECT 114.205 117.915 114.375 118.085 ;
        RECT 114.665 117.915 114.835 118.085 ;
        RECT 115.125 117.915 115.295 118.085 ;
        RECT 115.585 117.915 115.755 118.085 ;
        RECT 116.045 117.915 116.215 118.085 ;
        RECT 116.505 117.915 116.675 118.085 ;
        RECT 116.965 117.915 117.135 118.085 ;
        RECT 117.425 117.915 117.595 118.085 ;
        RECT 117.885 117.915 118.055 118.085 ;
        RECT 118.345 117.915 118.515 118.085 ;
        RECT 118.805 117.915 118.975 118.085 ;
        RECT 119.265 117.915 119.435 118.085 ;
        RECT 119.725 117.915 119.895 118.085 ;
        RECT 120.185 117.915 120.355 118.085 ;
        RECT 120.645 117.915 120.815 118.085 ;
        RECT 121.105 117.915 121.275 118.085 ;
        RECT 121.565 117.915 121.735 118.085 ;
        RECT 122.025 117.915 122.195 118.085 ;
        RECT 122.485 117.915 122.655 118.085 ;
        RECT 122.945 117.915 123.115 118.085 ;
        RECT 123.405 117.915 123.575 118.085 ;
        RECT 123.865 117.915 124.035 118.085 ;
        RECT 124.325 117.915 124.495 118.085 ;
        RECT 124.785 117.915 124.955 118.085 ;
        RECT 125.245 117.915 125.415 118.085 ;
        RECT 125.705 117.915 125.875 118.085 ;
        RECT 126.165 117.915 126.335 118.085 ;
        RECT 126.625 117.915 126.795 118.085 ;
        RECT 127.085 117.915 127.255 118.085 ;
        RECT 127.545 117.915 127.715 118.085 ;
        RECT 128.005 117.915 128.175 118.085 ;
        RECT 128.465 117.915 128.635 118.085 ;
        RECT 128.925 117.915 129.095 118.085 ;
        RECT 129.385 117.915 129.555 118.085 ;
        RECT 129.845 117.915 130.015 118.085 ;
        RECT 130.305 117.915 130.475 118.085 ;
        RECT 130.765 117.915 130.935 118.085 ;
        RECT 131.225 117.915 131.395 118.085 ;
        RECT 131.685 117.915 131.855 118.085 ;
        RECT 132.145 117.915 132.315 118.085 ;
        RECT 132.605 117.915 132.775 118.085 ;
        RECT 133.065 117.915 133.235 118.085 ;
        RECT 133.525 117.915 133.695 118.085 ;
        RECT 133.985 117.915 134.155 118.085 ;
        RECT 45.665 112.475 45.835 112.645 ;
        RECT 46.125 112.475 46.295 112.645 ;
        RECT 46.585 112.475 46.755 112.645 ;
        RECT 47.045 112.475 47.215 112.645 ;
        RECT 47.505 112.475 47.675 112.645 ;
        RECT 47.965 112.475 48.135 112.645 ;
        RECT 48.425 112.475 48.595 112.645 ;
        RECT 48.885 112.475 49.055 112.645 ;
        RECT 49.345 112.475 49.515 112.645 ;
        RECT 49.805 112.475 49.975 112.645 ;
        RECT 50.265 112.475 50.435 112.645 ;
        RECT 50.725 112.475 50.895 112.645 ;
        RECT 51.185 112.475 51.355 112.645 ;
        RECT 51.645 112.475 51.815 112.645 ;
        RECT 52.105 112.475 52.275 112.645 ;
        RECT 52.565 112.475 52.735 112.645 ;
        RECT 53.025 112.475 53.195 112.645 ;
        RECT 53.485 112.475 53.655 112.645 ;
        RECT 53.945 112.475 54.115 112.645 ;
        RECT 54.405 112.475 54.575 112.645 ;
        RECT 54.865 112.475 55.035 112.645 ;
        RECT 55.325 112.475 55.495 112.645 ;
        RECT 55.785 112.475 55.955 112.645 ;
        RECT 56.245 112.475 56.415 112.645 ;
        RECT 56.705 112.475 56.875 112.645 ;
        RECT 57.165 112.475 57.335 112.645 ;
        RECT 57.625 112.475 57.795 112.645 ;
        RECT 58.085 112.475 58.255 112.645 ;
        RECT 58.545 112.475 58.715 112.645 ;
        RECT 59.005 112.475 59.175 112.645 ;
        RECT 59.465 112.475 59.635 112.645 ;
        RECT 59.925 112.475 60.095 112.645 ;
        RECT 60.385 112.475 60.555 112.645 ;
        RECT 60.845 112.475 61.015 112.645 ;
        RECT 61.305 112.475 61.475 112.645 ;
        RECT 61.765 112.475 61.935 112.645 ;
        RECT 62.225 112.475 62.395 112.645 ;
        RECT 62.685 112.475 62.855 112.645 ;
        RECT 63.145 112.475 63.315 112.645 ;
        RECT 63.605 112.475 63.775 112.645 ;
        RECT 64.065 112.475 64.235 112.645 ;
        RECT 64.525 112.475 64.695 112.645 ;
        RECT 64.985 112.475 65.155 112.645 ;
        RECT 65.445 112.475 65.615 112.645 ;
        RECT 65.905 112.475 66.075 112.645 ;
        RECT 66.365 112.475 66.535 112.645 ;
        RECT 66.825 112.475 66.995 112.645 ;
        RECT 67.285 112.475 67.455 112.645 ;
        RECT 67.745 112.475 67.915 112.645 ;
        RECT 68.205 112.475 68.375 112.645 ;
        RECT 68.665 112.475 68.835 112.645 ;
        RECT 69.125 112.475 69.295 112.645 ;
        RECT 69.585 112.475 69.755 112.645 ;
        RECT 70.045 112.475 70.215 112.645 ;
        RECT 70.505 112.475 70.675 112.645 ;
        RECT 70.965 112.475 71.135 112.645 ;
        RECT 71.425 112.475 71.595 112.645 ;
        RECT 71.885 112.475 72.055 112.645 ;
        RECT 72.345 112.475 72.515 112.645 ;
        RECT 72.805 112.475 72.975 112.645 ;
        RECT 73.265 112.475 73.435 112.645 ;
        RECT 73.725 112.475 73.895 112.645 ;
        RECT 74.185 112.475 74.355 112.645 ;
        RECT 74.645 112.475 74.815 112.645 ;
        RECT 75.105 112.475 75.275 112.645 ;
        RECT 75.565 112.475 75.735 112.645 ;
        RECT 76.025 112.475 76.195 112.645 ;
        RECT 76.485 112.475 76.655 112.645 ;
        RECT 76.945 112.475 77.115 112.645 ;
        RECT 77.405 112.475 77.575 112.645 ;
        RECT 77.865 112.475 78.035 112.645 ;
        RECT 78.325 112.475 78.495 112.645 ;
        RECT 78.785 112.475 78.955 112.645 ;
        RECT 79.245 112.475 79.415 112.645 ;
        RECT 79.705 112.475 79.875 112.645 ;
        RECT 80.165 112.475 80.335 112.645 ;
        RECT 80.625 112.475 80.795 112.645 ;
        RECT 81.085 112.475 81.255 112.645 ;
        RECT 81.545 112.475 81.715 112.645 ;
        RECT 82.005 112.475 82.175 112.645 ;
        RECT 82.465 112.475 82.635 112.645 ;
        RECT 82.925 112.475 83.095 112.645 ;
        RECT 83.385 112.475 83.555 112.645 ;
        RECT 83.845 112.475 84.015 112.645 ;
        RECT 84.305 112.475 84.475 112.645 ;
        RECT 84.765 112.475 84.935 112.645 ;
        RECT 85.225 112.475 85.395 112.645 ;
        RECT 85.685 112.475 85.855 112.645 ;
        RECT 86.145 112.475 86.315 112.645 ;
        RECT 86.605 112.475 86.775 112.645 ;
        RECT 87.065 112.475 87.235 112.645 ;
        RECT 87.525 112.475 87.695 112.645 ;
        RECT 87.985 112.475 88.155 112.645 ;
        RECT 88.445 112.475 88.615 112.645 ;
        RECT 88.905 112.475 89.075 112.645 ;
        RECT 89.365 112.475 89.535 112.645 ;
        RECT 89.825 112.475 89.995 112.645 ;
        RECT 90.285 112.475 90.455 112.645 ;
        RECT 90.745 112.475 90.915 112.645 ;
        RECT 91.205 112.475 91.375 112.645 ;
        RECT 91.665 112.475 91.835 112.645 ;
        RECT 92.125 112.475 92.295 112.645 ;
        RECT 92.585 112.475 92.755 112.645 ;
        RECT 93.045 112.475 93.215 112.645 ;
        RECT 93.505 112.475 93.675 112.645 ;
        RECT 93.965 112.475 94.135 112.645 ;
        RECT 94.425 112.475 94.595 112.645 ;
        RECT 94.885 112.475 95.055 112.645 ;
        RECT 95.345 112.475 95.515 112.645 ;
        RECT 95.805 112.475 95.975 112.645 ;
        RECT 96.265 112.475 96.435 112.645 ;
        RECT 96.725 112.475 96.895 112.645 ;
        RECT 97.185 112.475 97.355 112.645 ;
        RECT 97.645 112.475 97.815 112.645 ;
        RECT 98.105 112.475 98.275 112.645 ;
        RECT 98.565 112.475 98.735 112.645 ;
        RECT 99.025 112.475 99.195 112.645 ;
        RECT 99.485 112.475 99.655 112.645 ;
        RECT 99.945 112.475 100.115 112.645 ;
        RECT 100.405 112.475 100.575 112.645 ;
        RECT 100.865 112.475 101.035 112.645 ;
        RECT 101.325 112.475 101.495 112.645 ;
        RECT 101.785 112.475 101.955 112.645 ;
        RECT 102.245 112.475 102.415 112.645 ;
        RECT 102.705 112.475 102.875 112.645 ;
        RECT 103.165 112.475 103.335 112.645 ;
        RECT 103.625 112.475 103.795 112.645 ;
        RECT 104.085 112.475 104.255 112.645 ;
        RECT 104.545 112.475 104.715 112.645 ;
        RECT 105.005 112.475 105.175 112.645 ;
        RECT 105.465 112.475 105.635 112.645 ;
        RECT 105.925 112.475 106.095 112.645 ;
        RECT 106.385 112.475 106.555 112.645 ;
        RECT 106.845 112.475 107.015 112.645 ;
        RECT 107.305 112.475 107.475 112.645 ;
        RECT 107.765 112.475 107.935 112.645 ;
        RECT 108.225 112.475 108.395 112.645 ;
        RECT 108.685 112.475 108.855 112.645 ;
        RECT 109.145 112.475 109.315 112.645 ;
        RECT 109.605 112.475 109.775 112.645 ;
        RECT 110.065 112.475 110.235 112.645 ;
        RECT 110.525 112.475 110.695 112.645 ;
        RECT 110.985 112.475 111.155 112.645 ;
        RECT 111.445 112.475 111.615 112.645 ;
        RECT 111.905 112.475 112.075 112.645 ;
        RECT 112.365 112.475 112.535 112.645 ;
        RECT 112.825 112.475 112.995 112.645 ;
        RECT 113.285 112.475 113.455 112.645 ;
        RECT 113.745 112.475 113.915 112.645 ;
        RECT 114.205 112.475 114.375 112.645 ;
        RECT 114.665 112.475 114.835 112.645 ;
        RECT 115.125 112.475 115.295 112.645 ;
        RECT 115.585 112.475 115.755 112.645 ;
        RECT 116.045 112.475 116.215 112.645 ;
        RECT 116.505 112.475 116.675 112.645 ;
        RECT 116.965 112.475 117.135 112.645 ;
        RECT 117.425 112.475 117.595 112.645 ;
        RECT 117.885 112.475 118.055 112.645 ;
        RECT 118.345 112.475 118.515 112.645 ;
        RECT 118.805 112.475 118.975 112.645 ;
        RECT 119.265 112.475 119.435 112.645 ;
        RECT 119.725 112.475 119.895 112.645 ;
        RECT 120.185 112.475 120.355 112.645 ;
        RECT 120.645 112.475 120.815 112.645 ;
        RECT 121.105 112.475 121.275 112.645 ;
        RECT 121.565 112.475 121.735 112.645 ;
        RECT 122.025 112.475 122.195 112.645 ;
        RECT 122.485 112.475 122.655 112.645 ;
        RECT 122.945 112.475 123.115 112.645 ;
        RECT 123.405 112.475 123.575 112.645 ;
        RECT 123.865 112.475 124.035 112.645 ;
        RECT 124.325 112.475 124.495 112.645 ;
        RECT 124.785 112.475 124.955 112.645 ;
        RECT 125.245 112.475 125.415 112.645 ;
        RECT 125.705 112.475 125.875 112.645 ;
        RECT 126.165 112.475 126.335 112.645 ;
        RECT 126.625 112.475 126.795 112.645 ;
        RECT 127.085 112.475 127.255 112.645 ;
        RECT 127.545 112.475 127.715 112.645 ;
        RECT 128.005 112.475 128.175 112.645 ;
        RECT 128.465 112.475 128.635 112.645 ;
        RECT 128.925 112.475 129.095 112.645 ;
        RECT 129.385 112.475 129.555 112.645 ;
        RECT 129.845 112.475 130.015 112.645 ;
        RECT 130.305 112.475 130.475 112.645 ;
        RECT 130.765 112.475 130.935 112.645 ;
        RECT 131.225 112.475 131.395 112.645 ;
        RECT 131.685 112.475 131.855 112.645 ;
        RECT 132.145 112.475 132.315 112.645 ;
        RECT 132.605 112.475 132.775 112.645 ;
        RECT 133.065 112.475 133.235 112.645 ;
        RECT 133.525 112.475 133.695 112.645 ;
        RECT 133.985 112.475 134.155 112.645 ;
        RECT 45.665 107.035 45.835 107.205 ;
        RECT 46.125 107.035 46.295 107.205 ;
        RECT 46.585 107.035 46.755 107.205 ;
        RECT 47.045 107.035 47.215 107.205 ;
        RECT 47.505 107.035 47.675 107.205 ;
        RECT 47.965 107.035 48.135 107.205 ;
        RECT 48.425 107.035 48.595 107.205 ;
        RECT 48.885 107.035 49.055 107.205 ;
        RECT 49.345 107.035 49.515 107.205 ;
        RECT 49.805 107.035 49.975 107.205 ;
        RECT 50.265 107.035 50.435 107.205 ;
        RECT 50.725 107.035 50.895 107.205 ;
        RECT 51.185 107.035 51.355 107.205 ;
        RECT 51.645 107.035 51.815 107.205 ;
        RECT 52.105 107.035 52.275 107.205 ;
        RECT 52.565 107.035 52.735 107.205 ;
        RECT 53.025 107.035 53.195 107.205 ;
        RECT 53.485 107.035 53.655 107.205 ;
        RECT 53.945 107.035 54.115 107.205 ;
        RECT 54.405 107.035 54.575 107.205 ;
        RECT 54.865 107.035 55.035 107.205 ;
        RECT 55.325 107.035 55.495 107.205 ;
        RECT 55.785 107.035 55.955 107.205 ;
        RECT 56.245 107.035 56.415 107.205 ;
        RECT 56.705 107.035 56.875 107.205 ;
        RECT 57.165 107.035 57.335 107.205 ;
        RECT 57.625 107.035 57.795 107.205 ;
        RECT 58.085 107.035 58.255 107.205 ;
        RECT 58.545 107.035 58.715 107.205 ;
        RECT 59.005 107.035 59.175 107.205 ;
        RECT 59.465 107.035 59.635 107.205 ;
        RECT 59.925 107.035 60.095 107.205 ;
        RECT 60.385 107.035 60.555 107.205 ;
        RECT 60.845 107.035 61.015 107.205 ;
        RECT 61.305 107.035 61.475 107.205 ;
        RECT 61.765 107.035 61.935 107.205 ;
        RECT 62.225 107.035 62.395 107.205 ;
        RECT 62.685 107.035 62.855 107.205 ;
        RECT 63.145 107.035 63.315 107.205 ;
        RECT 63.605 107.035 63.775 107.205 ;
        RECT 64.065 107.035 64.235 107.205 ;
        RECT 64.525 107.035 64.695 107.205 ;
        RECT 64.985 107.035 65.155 107.205 ;
        RECT 65.445 107.035 65.615 107.205 ;
        RECT 65.905 107.035 66.075 107.205 ;
        RECT 66.365 107.035 66.535 107.205 ;
        RECT 66.825 107.035 66.995 107.205 ;
        RECT 67.285 107.035 67.455 107.205 ;
        RECT 67.745 107.035 67.915 107.205 ;
        RECT 68.205 107.035 68.375 107.205 ;
        RECT 68.665 107.035 68.835 107.205 ;
        RECT 69.125 107.035 69.295 107.205 ;
        RECT 69.585 107.035 69.755 107.205 ;
        RECT 70.045 107.035 70.215 107.205 ;
        RECT 70.505 107.035 70.675 107.205 ;
        RECT 70.965 107.035 71.135 107.205 ;
        RECT 71.425 107.035 71.595 107.205 ;
        RECT 71.885 107.035 72.055 107.205 ;
        RECT 72.345 107.035 72.515 107.205 ;
        RECT 72.805 107.035 72.975 107.205 ;
        RECT 73.265 107.035 73.435 107.205 ;
        RECT 73.725 107.035 73.895 107.205 ;
        RECT 74.185 107.035 74.355 107.205 ;
        RECT 74.645 107.035 74.815 107.205 ;
        RECT 75.105 107.035 75.275 107.205 ;
        RECT 75.565 107.035 75.735 107.205 ;
        RECT 76.025 107.035 76.195 107.205 ;
        RECT 76.485 107.035 76.655 107.205 ;
        RECT 76.945 107.035 77.115 107.205 ;
        RECT 77.405 107.035 77.575 107.205 ;
        RECT 77.865 107.035 78.035 107.205 ;
        RECT 78.325 107.035 78.495 107.205 ;
        RECT 78.785 107.035 78.955 107.205 ;
        RECT 79.245 107.035 79.415 107.205 ;
        RECT 79.705 107.035 79.875 107.205 ;
        RECT 80.165 107.035 80.335 107.205 ;
        RECT 80.625 107.035 80.795 107.205 ;
        RECT 81.085 107.035 81.255 107.205 ;
        RECT 81.545 107.035 81.715 107.205 ;
        RECT 82.005 107.035 82.175 107.205 ;
        RECT 82.465 107.035 82.635 107.205 ;
        RECT 82.925 107.035 83.095 107.205 ;
        RECT 83.385 107.035 83.555 107.205 ;
        RECT 83.845 107.035 84.015 107.205 ;
        RECT 84.305 107.035 84.475 107.205 ;
        RECT 84.765 107.035 84.935 107.205 ;
        RECT 85.225 107.035 85.395 107.205 ;
        RECT 85.685 107.035 85.855 107.205 ;
        RECT 86.145 107.035 86.315 107.205 ;
        RECT 86.605 107.035 86.775 107.205 ;
        RECT 87.065 107.035 87.235 107.205 ;
        RECT 87.525 107.035 87.695 107.205 ;
        RECT 87.985 107.035 88.155 107.205 ;
        RECT 88.445 107.035 88.615 107.205 ;
        RECT 88.905 107.035 89.075 107.205 ;
        RECT 89.365 107.035 89.535 107.205 ;
        RECT 89.825 107.035 89.995 107.205 ;
        RECT 90.285 107.035 90.455 107.205 ;
        RECT 90.745 107.035 90.915 107.205 ;
        RECT 91.205 107.035 91.375 107.205 ;
        RECT 91.665 107.035 91.835 107.205 ;
        RECT 92.125 107.035 92.295 107.205 ;
        RECT 92.585 107.035 92.755 107.205 ;
        RECT 93.045 107.035 93.215 107.205 ;
        RECT 93.505 107.035 93.675 107.205 ;
        RECT 93.965 107.035 94.135 107.205 ;
        RECT 94.425 107.035 94.595 107.205 ;
        RECT 94.885 107.035 95.055 107.205 ;
        RECT 95.345 107.035 95.515 107.205 ;
        RECT 95.805 107.035 95.975 107.205 ;
        RECT 96.265 107.035 96.435 107.205 ;
        RECT 96.725 107.035 96.895 107.205 ;
        RECT 97.185 107.035 97.355 107.205 ;
        RECT 97.645 107.035 97.815 107.205 ;
        RECT 98.105 107.035 98.275 107.205 ;
        RECT 98.565 107.035 98.735 107.205 ;
        RECT 99.025 107.035 99.195 107.205 ;
        RECT 99.485 107.035 99.655 107.205 ;
        RECT 99.945 107.035 100.115 107.205 ;
        RECT 100.405 107.035 100.575 107.205 ;
        RECT 100.865 107.035 101.035 107.205 ;
        RECT 101.325 107.035 101.495 107.205 ;
        RECT 101.785 107.035 101.955 107.205 ;
        RECT 102.245 107.035 102.415 107.205 ;
        RECT 102.705 107.035 102.875 107.205 ;
        RECT 103.165 107.035 103.335 107.205 ;
        RECT 103.625 107.035 103.795 107.205 ;
        RECT 104.085 107.035 104.255 107.205 ;
        RECT 104.545 107.035 104.715 107.205 ;
        RECT 105.005 107.035 105.175 107.205 ;
        RECT 105.465 107.035 105.635 107.205 ;
        RECT 105.925 107.035 106.095 107.205 ;
        RECT 106.385 107.035 106.555 107.205 ;
        RECT 106.845 107.035 107.015 107.205 ;
        RECT 107.305 107.035 107.475 107.205 ;
        RECT 107.765 107.035 107.935 107.205 ;
        RECT 108.225 107.035 108.395 107.205 ;
        RECT 108.685 107.035 108.855 107.205 ;
        RECT 109.145 107.035 109.315 107.205 ;
        RECT 109.605 107.035 109.775 107.205 ;
        RECT 110.065 107.035 110.235 107.205 ;
        RECT 110.525 107.035 110.695 107.205 ;
        RECT 110.985 107.035 111.155 107.205 ;
        RECT 111.445 107.035 111.615 107.205 ;
        RECT 111.905 107.035 112.075 107.205 ;
        RECT 112.365 107.035 112.535 107.205 ;
        RECT 112.825 107.035 112.995 107.205 ;
        RECT 113.285 107.035 113.455 107.205 ;
        RECT 113.745 107.035 113.915 107.205 ;
        RECT 114.205 107.035 114.375 107.205 ;
        RECT 114.665 107.035 114.835 107.205 ;
        RECT 115.125 107.035 115.295 107.205 ;
        RECT 115.585 107.035 115.755 107.205 ;
        RECT 116.045 107.035 116.215 107.205 ;
        RECT 116.505 107.035 116.675 107.205 ;
        RECT 116.965 107.035 117.135 107.205 ;
        RECT 117.425 107.035 117.595 107.205 ;
        RECT 117.885 107.035 118.055 107.205 ;
        RECT 118.345 107.035 118.515 107.205 ;
        RECT 118.805 107.035 118.975 107.205 ;
        RECT 119.265 107.035 119.435 107.205 ;
        RECT 119.725 107.035 119.895 107.205 ;
        RECT 120.185 107.035 120.355 107.205 ;
        RECT 120.645 107.035 120.815 107.205 ;
        RECT 121.105 107.035 121.275 107.205 ;
        RECT 121.565 107.035 121.735 107.205 ;
        RECT 122.025 107.035 122.195 107.205 ;
        RECT 122.485 107.035 122.655 107.205 ;
        RECT 122.945 107.035 123.115 107.205 ;
        RECT 123.405 107.035 123.575 107.205 ;
        RECT 123.865 107.035 124.035 107.205 ;
        RECT 124.325 107.035 124.495 107.205 ;
        RECT 124.785 107.035 124.955 107.205 ;
        RECT 125.245 107.035 125.415 107.205 ;
        RECT 125.705 107.035 125.875 107.205 ;
        RECT 126.165 107.035 126.335 107.205 ;
        RECT 126.625 107.035 126.795 107.205 ;
        RECT 127.085 107.035 127.255 107.205 ;
        RECT 127.545 107.035 127.715 107.205 ;
        RECT 128.005 107.035 128.175 107.205 ;
        RECT 128.465 107.035 128.635 107.205 ;
        RECT 128.925 107.035 129.095 107.205 ;
        RECT 129.385 107.035 129.555 107.205 ;
        RECT 129.845 107.035 130.015 107.205 ;
        RECT 130.305 107.035 130.475 107.205 ;
        RECT 130.765 107.035 130.935 107.205 ;
        RECT 131.225 107.035 131.395 107.205 ;
        RECT 131.685 107.035 131.855 107.205 ;
        RECT 132.145 107.035 132.315 107.205 ;
        RECT 132.605 107.035 132.775 107.205 ;
        RECT 133.065 107.035 133.235 107.205 ;
        RECT 133.525 107.035 133.695 107.205 ;
        RECT 133.985 107.035 134.155 107.205 ;
        RECT 45.665 101.595 45.835 101.765 ;
        RECT 46.125 101.595 46.295 101.765 ;
        RECT 46.585 101.595 46.755 101.765 ;
        RECT 47.045 101.595 47.215 101.765 ;
        RECT 47.505 101.595 47.675 101.765 ;
        RECT 47.965 101.595 48.135 101.765 ;
        RECT 48.425 101.595 48.595 101.765 ;
        RECT 48.885 101.595 49.055 101.765 ;
        RECT 49.345 101.595 49.515 101.765 ;
        RECT 49.805 101.595 49.975 101.765 ;
        RECT 50.265 101.595 50.435 101.765 ;
        RECT 50.725 101.595 50.895 101.765 ;
        RECT 51.185 101.595 51.355 101.765 ;
        RECT 51.645 101.595 51.815 101.765 ;
        RECT 52.105 101.595 52.275 101.765 ;
        RECT 52.565 101.595 52.735 101.765 ;
        RECT 53.025 101.595 53.195 101.765 ;
        RECT 53.485 101.595 53.655 101.765 ;
        RECT 53.945 101.595 54.115 101.765 ;
        RECT 54.405 101.595 54.575 101.765 ;
        RECT 54.865 101.595 55.035 101.765 ;
        RECT 55.325 101.595 55.495 101.765 ;
        RECT 55.785 101.595 55.955 101.765 ;
        RECT 56.245 101.595 56.415 101.765 ;
        RECT 56.705 101.595 56.875 101.765 ;
        RECT 57.165 101.595 57.335 101.765 ;
        RECT 57.625 101.595 57.795 101.765 ;
        RECT 58.085 101.595 58.255 101.765 ;
        RECT 58.545 101.595 58.715 101.765 ;
        RECT 59.005 101.595 59.175 101.765 ;
        RECT 59.465 101.595 59.635 101.765 ;
        RECT 59.925 101.595 60.095 101.765 ;
        RECT 60.385 101.595 60.555 101.765 ;
        RECT 60.845 101.595 61.015 101.765 ;
        RECT 61.305 101.595 61.475 101.765 ;
        RECT 61.765 101.595 61.935 101.765 ;
        RECT 62.225 101.595 62.395 101.765 ;
        RECT 62.685 101.595 62.855 101.765 ;
        RECT 63.145 101.595 63.315 101.765 ;
        RECT 63.605 101.595 63.775 101.765 ;
        RECT 64.065 101.595 64.235 101.765 ;
        RECT 64.525 101.595 64.695 101.765 ;
        RECT 64.985 101.595 65.155 101.765 ;
        RECT 65.445 101.595 65.615 101.765 ;
        RECT 65.905 101.595 66.075 101.765 ;
        RECT 66.365 101.595 66.535 101.765 ;
        RECT 66.825 101.595 66.995 101.765 ;
        RECT 67.285 101.595 67.455 101.765 ;
        RECT 67.745 101.595 67.915 101.765 ;
        RECT 68.205 101.595 68.375 101.765 ;
        RECT 68.665 101.595 68.835 101.765 ;
        RECT 69.125 101.595 69.295 101.765 ;
        RECT 69.585 101.595 69.755 101.765 ;
        RECT 70.045 101.595 70.215 101.765 ;
        RECT 70.505 101.595 70.675 101.765 ;
        RECT 70.965 101.595 71.135 101.765 ;
        RECT 71.425 101.595 71.595 101.765 ;
        RECT 71.885 101.595 72.055 101.765 ;
        RECT 72.345 101.595 72.515 101.765 ;
        RECT 72.805 101.595 72.975 101.765 ;
        RECT 73.265 101.595 73.435 101.765 ;
        RECT 73.725 101.595 73.895 101.765 ;
        RECT 74.185 101.595 74.355 101.765 ;
        RECT 74.645 101.595 74.815 101.765 ;
        RECT 75.105 101.595 75.275 101.765 ;
        RECT 75.565 101.595 75.735 101.765 ;
        RECT 76.025 101.595 76.195 101.765 ;
        RECT 76.485 101.595 76.655 101.765 ;
        RECT 76.945 101.595 77.115 101.765 ;
        RECT 77.405 101.595 77.575 101.765 ;
        RECT 77.865 101.595 78.035 101.765 ;
        RECT 78.325 101.595 78.495 101.765 ;
        RECT 78.785 101.595 78.955 101.765 ;
        RECT 79.245 101.595 79.415 101.765 ;
        RECT 79.705 101.595 79.875 101.765 ;
        RECT 80.165 101.595 80.335 101.765 ;
        RECT 80.625 101.595 80.795 101.765 ;
        RECT 81.085 101.595 81.255 101.765 ;
        RECT 81.545 101.595 81.715 101.765 ;
        RECT 82.005 101.595 82.175 101.765 ;
        RECT 82.465 101.595 82.635 101.765 ;
        RECT 82.925 101.595 83.095 101.765 ;
        RECT 83.385 101.595 83.555 101.765 ;
        RECT 83.845 101.595 84.015 101.765 ;
        RECT 84.305 101.595 84.475 101.765 ;
        RECT 84.765 101.595 84.935 101.765 ;
        RECT 85.225 101.595 85.395 101.765 ;
        RECT 85.685 101.595 85.855 101.765 ;
        RECT 86.145 101.595 86.315 101.765 ;
        RECT 86.605 101.595 86.775 101.765 ;
        RECT 87.065 101.595 87.235 101.765 ;
        RECT 87.525 101.595 87.695 101.765 ;
        RECT 87.985 101.595 88.155 101.765 ;
        RECT 88.445 101.595 88.615 101.765 ;
        RECT 88.905 101.595 89.075 101.765 ;
        RECT 89.365 101.595 89.535 101.765 ;
        RECT 89.825 101.595 89.995 101.765 ;
        RECT 90.285 101.595 90.455 101.765 ;
        RECT 90.745 101.595 90.915 101.765 ;
        RECT 91.205 101.595 91.375 101.765 ;
        RECT 91.665 101.595 91.835 101.765 ;
        RECT 92.125 101.595 92.295 101.765 ;
        RECT 92.585 101.595 92.755 101.765 ;
        RECT 93.045 101.595 93.215 101.765 ;
        RECT 93.505 101.595 93.675 101.765 ;
        RECT 93.965 101.595 94.135 101.765 ;
        RECT 94.425 101.595 94.595 101.765 ;
        RECT 94.885 101.595 95.055 101.765 ;
        RECT 95.345 101.595 95.515 101.765 ;
        RECT 95.805 101.595 95.975 101.765 ;
        RECT 96.265 101.595 96.435 101.765 ;
        RECT 96.725 101.595 96.895 101.765 ;
        RECT 97.185 101.595 97.355 101.765 ;
        RECT 97.645 101.595 97.815 101.765 ;
        RECT 98.105 101.595 98.275 101.765 ;
        RECT 98.565 101.595 98.735 101.765 ;
        RECT 99.025 101.595 99.195 101.765 ;
        RECT 99.485 101.595 99.655 101.765 ;
        RECT 99.945 101.595 100.115 101.765 ;
        RECT 100.405 101.595 100.575 101.765 ;
        RECT 100.865 101.595 101.035 101.765 ;
        RECT 101.325 101.595 101.495 101.765 ;
        RECT 101.785 101.595 101.955 101.765 ;
        RECT 102.245 101.595 102.415 101.765 ;
        RECT 102.705 101.595 102.875 101.765 ;
        RECT 103.165 101.595 103.335 101.765 ;
        RECT 103.625 101.595 103.795 101.765 ;
        RECT 104.085 101.595 104.255 101.765 ;
        RECT 104.545 101.595 104.715 101.765 ;
        RECT 105.005 101.595 105.175 101.765 ;
        RECT 105.465 101.595 105.635 101.765 ;
        RECT 105.925 101.595 106.095 101.765 ;
        RECT 106.385 101.595 106.555 101.765 ;
        RECT 106.845 101.595 107.015 101.765 ;
        RECT 107.305 101.595 107.475 101.765 ;
        RECT 107.765 101.595 107.935 101.765 ;
        RECT 108.225 101.595 108.395 101.765 ;
        RECT 108.685 101.595 108.855 101.765 ;
        RECT 109.145 101.595 109.315 101.765 ;
        RECT 109.605 101.595 109.775 101.765 ;
        RECT 110.065 101.595 110.235 101.765 ;
        RECT 110.525 101.595 110.695 101.765 ;
        RECT 110.985 101.595 111.155 101.765 ;
        RECT 111.445 101.595 111.615 101.765 ;
        RECT 111.905 101.595 112.075 101.765 ;
        RECT 112.365 101.595 112.535 101.765 ;
        RECT 112.825 101.595 112.995 101.765 ;
        RECT 113.285 101.595 113.455 101.765 ;
        RECT 113.745 101.595 113.915 101.765 ;
        RECT 114.205 101.595 114.375 101.765 ;
        RECT 114.665 101.595 114.835 101.765 ;
        RECT 115.125 101.595 115.295 101.765 ;
        RECT 115.585 101.595 115.755 101.765 ;
        RECT 116.045 101.595 116.215 101.765 ;
        RECT 116.505 101.595 116.675 101.765 ;
        RECT 116.965 101.595 117.135 101.765 ;
        RECT 117.425 101.595 117.595 101.765 ;
        RECT 117.885 101.595 118.055 101.765 ;
        RECT 118.345 101.595 118.515 101.765 ;
        RECT 118.805 101.595 118.975 101.765 ;
        RECT 119.265 101.595 119.435 101.765 ;
        RECT 119.725 101.595 119.895 101.765 ;
        RECT 120.185 101.595 120.355 101.765 ;
        RECT 120.645 101.595 120.815 101.765 ;
        RECT 121.105 101.595 121.275 101.765 ;
        RECT 121.565 101.595 121.735 101.765 ;
        RECT 122.025 101.595 122.195 101.765 ;
        RECT 122.485 101.595 122.655 101.765 ;
        RECT 122.945 101.595 123.115 101.765 ;
        RECT 123.405 101.595 123.575 101.765 ;
        RECT 123.865 101.595 124.035 101.765 ;
        RECT 124.325 101.595 124.495 101.765 ;
        RECT 124.785 101.595 124.955 101.765 ;
        RECT 125.245 101.595 125.415 101.765 ;
        RECT 125.705 101.595 125.875 101.765 ;
        RECT 126.165 101.595 126.335 101.765 ;
        RECT 126.625 101.595 126.795 101.765 ;
        RECT 127.085 101.595 127.255 101.765 ;
        RECT 127.545 101.595 127.715 101.765 ;
        RECT 128.005 101.595 128.175 101.765 ;
        RECT 128.465 101.595 128.635 101.765 ;
        RECT 128.925 101.595 129.095 101.765 ;
        RECT 129.385 101.595 129.555 101.765 ;
        RECT 129.845 101.595 130.015 101.765 ;
        RECT 130.305 101.595 130.475 101.765 ;
        RECT 130.765 101.595 130.935 101.765 ;
        RECT 131.225 101.595 131.395 101.765 ;
        RECT 131.685 101.595 131.855 101.765 ;
        RECT 132.145 101.595 132.315 101.765 ;
        RECT 132.605 101.595 132.775 101.765 ;
        RECT 133.065 101.595 133.235 101.765 ;
        RECT 133.525 101.595 133.695 101.765 ;
        RECT 133.985 101.595 134.155 101.765 ;
        RECT 45.665 96.155 45.835 96.325 ;
        RECT 46.125 96.155 46.295 96.325 ;
        RECT 46.585 96.155 46.755 96.325 ;
        RECT 47.045 96.155 47.215 96.325 ;
        RECT 47.505 96.155 47.675 96.325 ;
        RECT 47.965 96.155 48.135 96.325 ;
        RECT 48.425 96.155 48.595 96.325 ;
        RECT 48.885 96.155 49.055 96.325 ;
        RECT 49.345 96.155 49.515 96.325 ;
        RECT 49.805 96.155 49.975 96.325 ;
        RECT 50.265 96.155 50.435 96.325 ;
        RECT 50.725 96.155 50.895 96.325 ;
        RECT 51.185 96.155 51.355 96.325 ;
        RECT 51.645 96.155 51.815 96.325 ;
        RECT 52.105 96.155 52.275 96.325 ;
        RECT 52.565 96.155 52.735 96.325 ;
        RECT 53.025 96.155 53.195 96.325 ;
        RECT 53.485 96.155 53.655 96.325 ;
        RECT 53.945 96.155 54.115 96.325 ;
        RECT 54.405 96.155 54.575 96.325 ;
        RECT 54.865 96.155 55.035 96.325 ;
        RECT 55.325 96.155 55.495 96.325 ;
        RECT 55.785 96.155 55.955 96.325 ;
        RECT 56.245 96.155 56.415 96.325 ;
        RECT 56.705 96.155 56.875 96.325 ;
        RECT 57.165 96.155 57.335 96.325 ;
        RECT 57.625 96.155 57.795 96.325 ;
        RECT 58.085 96.155 58.255 96.325 ;
        RECT 58.545 96.155 58.715 96.325 ;
        RECT 59.005 96.155 59.175 96.325 ;
        RECT 59.465 96.155 59.635 96.325 ;
        RECT 59.925 96.155 60.095 96.325 ;
        RECT 60.385 96.155 60.555 96.325 ;
        RECT 60.845 96.155 61.015 96.325 ;
        RECT 61.305 96.155 61.475 96.325 ;
        RECT 61.765 96.155 61.935 96.325 ;
        RECT 62.225 96.155 62.395 96.325 ;
        RECT 62.685 96.155 62.855 96.325 ;
        RECT 63.145 96.155 63.315 96.325 ;
        RECT 63.605 96.155 63.775 96.325 ;
        RECT 64.065 96.155 64.235 96.325 ;
        RECT 64.525 96.155 64.695 96.325 ;
        RECT 64.985 96.155 65.155 96.325 ;
        RECT 65.445 96.155 65.615 96.325 ;
        RECT 65.905 96.155 66.075 96.325 ;
        RECT 66.365 96.155 66.535 96.325 ;
        RECT 66.825 96.155 66.995 96.325 ;
        RECT 67.285 96.155 67.455 96.325 ;
        RECT 67.745 96.155 67.915 96.325 ;
        RECT 68.205 96.155 68.375 96.325 ;
        RECT 68.665 96.155 68.835 96.325 ;
        RECT 69.125 96.155 69.295 96.325 ;
        RECT 69.585 96.155 69.755 96.325 ;
        RECT 70.045 96.155 70.215 96.325 ;
        RECT 70.505 96.155 70.675 96.325 ;
        RECT 70.965 96.155 71.135 96.325 ;
        RECT 71.425 96.155 71.595 96.325 ;
        RECT 71.885 96.155 72.055 96.325 ;
        RECT 72.345 96.155 72.515 96.325 ;
        RECT 72.805 96.155 72.975 96.325 ;
        RECT 73.265 96.155 73.435 96.325 ;
        RECT 73.725 96.155 73.895 96.325 ;
        RECT 74.185 96.155 74.355 96.325 ;
        RECT 74.645 96.155 74.815 96.325 ;
        RECT 75.105 96.155 75.275 96.325 ;
        RECT 75.565 96.155 75.735 96.325 ;
        RECT 76.025 96.155 76.195 96.325 ;
        RECT 76.485 96.155 76.655 96.325 ;
        RECT 76.945 96.155 77.115 96.325 ;
        RECT 77.405 96.155 77.575 96.325 ;
        RECT 77.865 96.155 78.035 96.325 ;
        RECT 78.325 96.155 78.495 96.325 ;
        RECT 78.785 96.155 78.955 96.325 ;
        RECT 79.245 96.155 79.415 96.325 ;
        RECT 79.705 96.155 79.875 96.325 ;
        RECT 80.165 96.155 80.335 96.325 ;
        RECT 80.625 96.155 80.795 96.325 ;
        RECT 81.085 96.155 81.255 96.325 ;
        RECT 81.545 96.155 81.715 96.325 ;
        RECT 82.005 96.155 82.175 96.325 ;
        RECT 82.465 96.155 82.635 96.325 ;
        RECT 82.925 96.155 83.095 96.325 ;
        RECT 83.385 96.155 83.555 96.325 ;
        RECT 83.845 96.155 84.015 96.325 ;
        RECT 84.305 96.155 84.475 96.325 ;
        RECT 84.765 96.155 84.935 96.325 ;
        RECT 85.225 96.155 85.395 96.325 ;
        RECT 85.685 96.155 85.855 96.325 ;
        RECT 86.145 96.155 86.315 96.325 ;
        RECT 86.605 96.155 86.775 96.325 ;
        RECT 87.065 96.155 87.235 96.325 ;
        RECT 87.525 96.155 87.695 96.325 ;
        RECT 87.985 96.155 88.155 96.325 ;
        RECT 88.445 96.155 88.615 96.325 ;
        RECT 88.905 96.155 89.075 96.325 ;
        RECT 89.365 96.155 89.535 96.325 ;
        RECT 89.825 96.155 89.995 96.325 ;
        RECT 90.285 96.155 90.455 96.325 ;
        RECT 90.745 96.155 90.915 96.325 ;
        RECT 91.205 96.155 91.375 96.325 ;
        RECT 91.665 96.155 91.835 96.325 ;
        RECT 92.125 96.155 92.295 96.325 ;
        RECT 92.585 96.155 92.755 96.325 ;
        RECT 93.045 96.155 93.215 96.325 ;
        RECT 93.505 96.155 93.675 96.325 ;
        RECT 93.965 96.155 94.135 96.325 ;
        RECT 94.425 96.155 94.595 96.325 ;
        RECT 94.885 96.155 95.055 96.325 ;
        RECT 95.345 96.155 95.515 96.325 ;
        RECT 95.805 96.155 95.975 96.325 ;
        RECT 96.265 96.155 96.435 96.325 ;
        RECT 96.725 96.155 96.895 96.325 ;
        RECT 97.185 96.155 97.355 96.325 ;
        RECT 97.645 96.155 97.815 96.325 ;
        RECT 98.105 96.155 98.275 96.325 ;
        RECT 98.565 96.155 98.735 96.325 ;
        RECT 99.025 96.155 99.195 96.325 ;
        RECT 99.485 96.155 99.655 96.325 ;
        RECT 99.945 96.155 100.115 96.325 ;
        RECT 100.405 96.155 100.575 96.325 ;
        RECT 100.865 96.155 101.035 96.325 ;
        RECT 101.325 96.155 101.495 96.325 ;
        RECT 101.785 96.155 101.955 96.325 ;
        RECT 102.245 96.155 102.415 96.325 ;
        RECT 102.705 96.155 102.875 96.325 ;
        RECT 103.165 96.155 103.335 96.325 ;
        RECT 103.625 96.155 103.795 96.325 ;
        RECT 104.085 96.155 104.255 96.325 ;
        RECT 104.545 96.155 104.715 96.325 ;
        RECT 105.005 96.155 105.175 96.325 ;
        RECT 105.465 96.155 105.635 96.325 ;
        RECT 105.925 96.155 106.095 96.325 ;
        RECT 106.385 96.155 106.555 96.325 ;
        RECT 106.845 96.155 107.015 96.325 ;
        RECT 107.305 96.155 107.475 96.325 ;
        RECT 107.765 96.155 107.935 96.325 ;
        RECT 108.225 96.155 108.395 96.325 ;
        RECT 108.685 96.155 108.855 96.325 ;
        RECT 109.145 96.155 109.315 96.325 ;
        RECT 109.605 96.155 109.775 96.325 ;
        RECT 110.065 96.155 110.235 96.325 ;
        RECT 110.525 96.155 110.695 96.325 ;
        RECT 110.985 96.155 111.155 96.325 ;
        RECT 111.445 96.155 111.615 96.325 ;
        RECT 111.905 96.155 112.075 96.325 ;
        RECT 112.365 96.155 112.535 96.325 ;
        RECT 112.825 96.155 112.995 96.325 ;
        RECT 113.285 96.155 113.455 96.325 ;
        RECT 113.745 96.155 113.915 96.325 ;
        RECT 114.205 96.155 114.375 96.325 ;
        RECT 114.665 96.155 114.835 96.325 ;
        RECT 115.125 96.155 115.295 96.325 ;
        RECT 115.585 96.155 115.755 96.325 ;
        RECT 116.045 96.155 116.215 96.325 ;
        RECT 116.505 96.155 116.675 96.325 ;
        RECT 116.965 96.155 117.135 96.325 ;
        RECT 117.425 96.155 117.595 96.325 ;
        RECT 117.885 96.155 118.055 96.325 ;
        RECT 118.345 96.155 118.515 96.325 ;
        RECT 118.805 96.155 118.975 96.325 ;
        RECT 119.265 96.155 119.435 96.325 ;
        RECT 119.725 96.155 119.895 96.325 ;
        RECT 120.185 96.155 120.355 96.325 ;
        RECT 120.645 96.155 120.815 96.325 ;
        RECT 121.105 96.155 121.275 96.325 ;
        RECT 121.565 96.155 121.735 96.325 ;
        RECT 122.025 96.155 122.195 96.325 ;
        RECT 122.485 96.155 122.655 96.325 ;
        RECT 122.945 96.155 123.115 96.325 ;
        RECT 123.405 96.155 123.575 96.325 ;
        RECT 123.865 96.155 124.035 96.325 ;
        RECT 124.325 96.155 124.495 96.325 ;
        RECT 124.785 96.155 124.955 96.325 ;
        RECT 125.245 96.155 125.415 96.325 ;
        RECT 125.705 96.155 125.875 96.325 ;
        RECT 126.165 96.155 126.335 96.325 ;
        RECT 126.625 96.155 126.795 96.325 ;
        RECT 127.085 96.155 127.255 96.325 ;
        RECT 127.545 96.155 127.715 96.325 ;
        RECT 128.005 96.155 128.175 96.325 ;
        RECT 128.465 96.155 128.635 96.325 ;
        RECT 128.925 96.155 129.095 96.325 ;
        RECT 129.385 96.155 129.555 96.325 ;
        RECT 129.845 96.155 130.015 96.325 ;
        RECT 130.305 96.155 130.475 96.325 ;
        RECT 130.765 96.155 130.935 96.325 ;
        RECT 131.225 96.155 131.395 96.325 ;
        RECT 131.685 96.155 131.855 96.325 ;
        RECT 132.145 96.155 132.315 96.325 ;
        RECT 132.605 96.155 132.775 96.325 ;
        RECT 133.065 96.155 133.235 96.325 ;
        RECT 133.525 96.155 133.695 96.325 ;
        RECT 133.985 96.155 134.155 96.325 ;
        RECT 45.665 90.715 45.835 90.885 ;
        RECT 46.125 90.715 46.295 90.885 ;
        RECT 46.585 90.715 46.755 90.885 ;
        RECT 47.045 90.715 47.215 90.885 ;
        RECT 47.505 90.715 47.675 90.885 ;
        RECT 47.965 90.715 48.135 90.885 ;
        RECT 48.425 90.715 48.595 90.885 ;
        RECT 48.885 90.715 49.055 90.885 ;
        RECT 49.345 90.715 49.515 90.885 ;
        RECT 49.805 90.715 49.975 90.885 ;
        RECT 50.265 90.715 50.435 90.885 ;
        RECT 50.725 90.715 50.895 90.885 ;
        RECT 51.185 90.715 51.355 90.885 ;
        RECT 51.645 90.715 51.815 90.885 ;
        RECT 52.105 90.715 52.275 90.885 ;
        RECT 52.565 90.715 52.735 90.885 ;
        RECT 53.025 90.715 53.195 90.885 ;
        RECT 53.485 90.715 53.655 90.885 ;
        RECT 53.945 90.715 54.115 90.885 ;
        RECT 54.405 90.715 54.575 90.885 ;
        RECT 54.865 90.715 55.035 90.885 ;
        RECT 55.325 90.715 55.495 90.885 ;
        RECT 55.785 90.715 55.955 90.885 ;
        RECT 56.245 90.715 56.415 90.885 ;
        RECT 56.705 90.715 56.875 90.885 ;
        RECT 57.165 90.715 57.335 90.885 ;
        RECT 57.625 90.715 57.795 90.885 ;
        RECT 58.085 90.715 58.255 90.885 ;
        RECT 58.545 90.715 58.715 90.885 ;
        RECT 59.005 90.715 59.175 90.885 ;
        RECT 59.465 90.715 59.635 90.885 ;
        RECT 59.925 90.715 60.095 90.885 ;
        RECT 60.385 90.715 60.555 90.885 ;
        RECT 60.845 90.715 61.015 90.885 ;
        RECT 61.305 90.715 61.475 90.885 ;
        RECT 61.765 90.715 61.935 90.885 ;
        RECT 62.225 90.715 62.395 90.885 ;
        RECT 62.685 90.715 62.855 90.885 ;
        RECT 63.145 90.715 63.315 90.885 ;
        RECT 63.605 90.715 63.775 90.885 ;
        RECT 64.065 90.715 64.235 90.885 ;
        RECT 64.525 90.715 64.695 90.885 ;
        RECT 64.985 90.715 65.155 90.885 ;
        RECT 65.445 90.715 65.615 90.885 ;
        RECT 65.905 90.715 66.075 90.885 ;
        RECT 66.365 90.715 66.535 90.885 ;
        RECT 66.825 90.715 66.995 90.885 ;
        RECT 67.285 90.715 67.455 90.885 ;
        RECT 67.745 90.715 67.915 90.885 ;
        RECT 68.205 90.715 68.375 90.885 ;
        RECT 68.665 90.715 68.835 90.885 ;
        RECT 69.125 90.715 69.295 90.885 ;
        RECT 69.585 90.715 69.755 90.885 ;
        RECT 70.045 90.715 70.215 90.885 ;
        RECT 70.505 90.715 70.675 90.885 ;
        RECT 70.965 90.715 71.135 90.885 ;
        RECT 71.425 90.715 71.595 90.885 ;
        RECT 71.885 90.715 72.055 90.885 ;
        RECT 72.345 90.715 72.515 90.885 ;
        RECT 72.805 90.715 72.975 90.885 ;
        RECT 73.265 90.715 73.435 90.885 ;
        RECT 73.725 90.715 73.895 90.885 ;
        RECT 74.185 90.715 74.355 90.885 ;
        RECT 74.645 90.715 74.815 90.885 ;
        RECT 75.105 90.715 75.275 90.885 ;
        RECT 75.565 90.715 75.735 90.885 ;
        RECT 76.025 90.715 76.195 90.885 ;
        RECT 76.485 90.715 76.655 90.885 ;
        RECT 76.945 90.715 77.115 90.885 ;
        RECT 77.405 90.715 77.575 90.885 ;
        RECT 77.865 90.715 78.035 90.885 ;
        RECT 78.325 90.715 78.495 90.885 ;
        RECT 78.785 90.715 78.955 90.885 ;
        RECT 79.245 90.715 79.415 90.885 ;
        RECT 79.705 90.715 79.875 90.885 ;
        RECT 80.165 90.715 80.335 90.885 ;
        RECT 80.625 90.715 80.795 90.885 ;
        RECT 81.085 90.715 81.255 90.885 ;
        RECT 81.545 90.715 81.715 90.885 ;
        RECT 82.005 90.715 82.175 90.885 ;
        RECT 82.465 90.715 82.635 90.885 ;
        RECT 82.925 90.715 83.095 90.885 ;
        RECT 83.385 90.715 83.555 90.885 ;
        RECT 83.845 90.715 84.015 90.885 ;
        RECT 84.305 90.715 84.475 90.885 ;
        RECT 84.765 90.715 84.935 90.885 ;
        RECT 85.225 90.715 85.395 90.885 ;
        RECT 85.685 90.715 85.855 90.885 ;
        RECT 86.145 90.715 86.315 90.885 ;
        RECT 86.605 90.715 86.775 90.885 ;
        RECT 87.065 90.715 87.235 90.885 ;
        RECT 87.525 90.715 87.695 90.885 ;
        RECT 87.985 90.715 88.155 90.885 ;
        RECT 88.445 90.715 88.615 90.885 ;
        RECT 88.905 90.715 89.075 90.885 ;
        RECT 89.365 90.715 89.535 90.885 ;
        RECT 89.825 90.715 89.995 90.885 ;
        RECT 90.285 90.715 90.455 90.885 ;
        RECT 90.745 90.715 90.915 90.885 ;
        RECT 91.205 90.715 91.375 90.885 ;
        RECT 91.665 90.715 91.835 90.885 ;
        RECT 92.125 90.715 92.295 90.885 ;
        RECT 92.585 90.715 92.755 90.885 ;
        RECT 93.045 90.715 93.215 90.885 ;
        RECT 93.505 90.715 93.675 90.885 ;
        RECT 93.965 90.715 94.135 90.885 ;
        RECT 94.425 90.715 94.595 90.885 ;
        RECT 94.885 90.715 95.055 90.885 ;
        RECT 95.345 90.715 95.515 90.885 ;
        RECT 95.805 90.715 95.975 90.885 ;
        RECT 96.265 90.715 96.435 90.885 ;
        RECT 96.725 90.715 96.895 90.885 ;
        RECT 97.185 90.715 97.355 90.885 ;
        RECT 97.645 90.715 97.815 90.885 ;
        RECT 98.105 90.715 98.275 90.885 ;
        RECT 98.565 90.715 98.735 90.885 ;
        RECT 99.025 90.715 99.195 90.885 ;
        RECT 99.485 90.715 99.655 90.885 ;
        RECT 99.945 90.715 100.115 90.885 ;
        RECT 100.405 90.715 100.575 90.885 ;
        RECT 100.865 90.715 101.035 90.885 ;
        RECT 101.325 90.715 101.495 90.885 ;
        RECT 101.785 90.715 101.955 90.885 ;
        RECT 102.245 90.715 102.415 90.885 ;
        RECT 102.705 90.715 102.875 90.885 ;
        RECT 103.165 90.715 103.335 90.885 ;
        RECT 103.625 90.715 103.795 90.885 ;
        RECT 104.085 90.715 104.255 90.885 ;
        RECT 104.545 90.715 104.715 90.885 ;
        RECT 105.005 90.715 105.175 90.885 ;
        RECT 105.465 90.715 105.635 90.885 ;
        RECT 105.925 90.715 106.095 90.885 ;
        RECT 106.385 90.715 106.555 90.885 ;
        RECT 106.845 90.715 107.015 90.885 ;
        RECT 107.305 90.715 107.475 90.885 ;
        RECT 107.765 90.715 107.935 90.885 ;
        RECT 108.225 90.715 108.395 90.885 ;
        RECT 108.685 90.715 108.855 90.885 ;
        RECT 109.145 90.715 109.315 90.885 ;
        RECT 109.605 90.715 109.775 90.885 ;
        RECT 110.065 90.715 110.235 90.885 ;
        RECT 110.525 90.715 110.695 90.885 ;
        RECT 110.985 90.715 111.155 90.885 ;
        RECT 111.445 90.715 111.615 90.885 ;
        RECT 111.905 90.715 112.075 90.885 ;
        RECT 112.365 90.715 112.535 90.885 ;
        RECT 112.825 90.715 112.995 90.885 ;
        RECT 113.285 90.715 113.455 90.885 ;
        RECT 113.745 90.715 113.915 90.885 ;
        RECT 114.205 90.715 114.375 90.885 ;
        RECT 114.665 90.715 114.835 90.885 ;
        RECT 115.125 90.715 115.295 90.885 ;
        RECT 115.585 90.715 115.755 90.885 ;
        RECT 116.045 90.715 116.215 90.885 ;
        RECT 116.505 90.715 116.675 90.885 ;
        RECT 116.965 90.715 117.135 90.885 ;
        RECT 117.425 90.715 117.595 90.885 ;
        RECT 117.885 90.715 118.055 90.885 ;
        RECT 118.345 90.715 118.515 90.885 ;
        RECT 118.805 90.715 118.975 90.885 ;
        RECT 119.265 90.715 119.435 90.885 ;
        RECT 119.725 90.715 119.895 90.885 ;
        RECT 120.185 90.715 120.355 90.885 ;
        RECT 120.645 90.715 120.815 90.885 ;
        RECT 121.105 90.715 121.275 90.885 ;
        RECT 121.565 90.715 121.735 90.885 ;
        RECT 122.025 90.715 122.195 90.885 ;
        RECT 122.485 90.715 122.655 90.885 ;
        RECT 122.945 90.715 123.115 90.885 ;
        RECT 123.405 90.715 123.575 90.885 ;
        RECT 123.865 90.715 124.035 90.885 ;
        RECT 124.325 90.715 124.495 90.885 ;
        RECT 124.785 90.715 124.955 90.885 ;
        RECT 125.245 90.715 125.415 90.885 ;
        RECT 125.705 90.715 125.875 90.885 ;
        RECT 126.165 90.715 126.335 90.885 ;
        RECT 126.625 90.715 126.795 90.885 ;
        RECT 127.085 90.715 127.255 90.885 ;
        RECT 127.545 90.715 127.715 90.885 ;
        RECT 128.005 90.715 128.175 90.885 ;
        RECT 128.465 90.715 128.635 90.885 ;
        RECT 128.925 90.715 129.095 90.885 ;
        RECT 129.385 90.715 129.555 90.885 ;
        RECT 129.845 90.715 130.015 90.885 ;
        RECT 130.305 90.715 130.475 90.885 ;
        RECT 130.765 90.715 130.935 90.885 ;
        RECT 131.225 90.715 131.395 90.885 ;
        RECT 131.685 90.715 131.855 90.885 ;
        RECT 132.145 90.715 132.315 90.885 ;
        RECT 132.605 90.715 132.775 90.885 ;
        RECT 133.065 90.715 133.235 90.885 ;
        RECT 133.525 90.715 133.695 90.885 ;
        RECT 133.985 90.715 134.155 90.885 ;
        RECT 45.665 85.275 45.835 85.445 ;
        RECT 46.125 85.275 46.295 85.445 ;
        RECT 46.585 85.275 46.755 85.445 ;
        RECT 47.045 85.275 47.215 85.445 ;
        RECT 47.505 85.275 47.675 85.445 ;
        RECT 47.965 85.275 48.135 85.445 ;
        RECT 48.425 85.275 48.595 85.445 ;
        RECT 48.885 85.275 49.055 85.445 ;
        RECT 49.345 85.275 49.515 85.445 ;
        RECT 49.805 85.275 49.975 85.445 ;
        RECT 50.265 85.275 50.435 85.445 ;
        RECT 50.725 85.275 50.895 85.445 ;
        RECT 51.185 85.275 51.355 85.445 ;
        RECT 51.645 85.275 51.815 85.445 ;
        RECT 52.105 85.275 52.275 85.445 ;
        RECT 52.565 85.275 52.735 85.445 ;
        RECT 53.025 85.275 53.195 85.445 ;
        RECT 53.485 85.275 53.655 85.445 ;
        RECT 53.945 85.275 54.115 85.445 ;
        RECT 54.405 85.275 54.575 85.445 ;
        RECT 54.865 85.275 55.035 85.445 ;
        RECT 55.325 85.275 55.495 85.445 ;
        RECT 55.785 85.275 55.955 85.445 ;
        RECT 56.245 85.275 56.415 85.445 ;
        RECT 56.705 85.275 56.875 85.445 ;
        RECT 57.165 85.275 57.335 85.445 ;
        RECT 57.625 85.275 57.795 85.445 ;
        RECT 58.085 85.275 58.255 85.445 ;
        RECT 58.545 85.275 58.715 85.445 ;
        RECT 59.005 85.275 59.175 85.445 ;
        RECT 59.465 85.275 59.635 85.445 ;
        RECT 59.925 85.275 60.095 85.445 ;
        RECT 60.385 85.275 60.555 85.445 ;
        RECT 60.845 85.275 61.015 85.445 ;
        RECT 61.305 85.275 61.475 85.445 ;
        RECT 61.765 85.275 61.935 85.445 ;
        RECT 62.225 85.275 62.395 85.445 ;
        RECT 62.685 85.275 62.855 85.445 ;
        RECT 63.145 85.275 63.315 85.445 ;
        RECT 63.605 85.275 63.775 85.445 ;
        RECT 64.065 85.275 64.235 85.445 ;
        RECT 64.525 85.275 64.695 85.445 ;
        RECT 64.985 85.275 65.155 85.445 ;
        RECT 65.445 85.275 65.615 85.445 ;
        RECT 65.905 85.275 66.075 85.445 ;
        RECT 66.365 85.275 66.535 85.445 ;
        RECT 66.825 85.275 66.995 85.445 ;
        RECT 67.285 85.275 67.455 85.445 ;
        RECT 67.745 85.275 67.915 85.445 ;
        RECT 68.205 85.275 68.375 85.445 ;
        RECT 68.665 85.275 68.835 85.445 ;
        RECT 69.125 85.275 69.295 85.445 ;
        RECT 69.585 85.275 69.755 85.445 ;
        RECT 70.045 85.275 70.215 85.445 ;
        RECT 70.505 85.275 70.675 85.445 ;
        RECT 70.965 85.275 71.135 85.445 ;
        RECT 71.425 85.275 71.595 85.445 ;
        RECT 71.885 85.275 72.055 85.445 ;
        RECT 72.345 85.275 72.515 85.445 ;
        RECT 72.805 85.275 72.975 85.445 ;
        RECT 73.265 85.275 73.435 85.445 ;
        RECT 73.725 85.275 73.895 85.445 ;
        RECT 74.185 85.275 74.355 85.445 ;
        RECT 74.645 85.275 74.815 85.445 ;
        RECT 75.105 85.275 75.275 85.445 ;
        RECT 75.565 85.275 75.735 85.445 ;
        RECT 76.025 85.275 76.195 85.445 ;
        RECT 76.485 85.275 76.655 85.445 ;
        RECT 76.945 85.275 77.115 85.445 ;
        RECT 77.405 85.275 77.575 85.445 ;
        RECT 77.865 85.275 78.035 85.445 ;
        RECT 78.325 85.275 78.495 85.445 ;
        RECT 78.785 85.275 78.955 85.445 ;
        RECT 79.245 85.275 79.415 85.445 ;
        RECT 79.705 85.275 79.875 85.445 ;
        RECT 80.165 85.275 80.335 85.445 ;
        RECT 80.625 85.275 80.795 85.445 ;
        RECT 81.085 85.275 81.255 85.445 ;
        RECT 81.545 85.275 81.715 85.445 ;
        RECT 82.005 85.275 82.175 85.445 ;
        RECT 82.465 85.275 82.635 85.445 ;
        RECT 82.925 85.275 83.095 85.445 ;
        RECT 83.385 85.275 83.555 85.445 ;
        RECT 83.845 85.275 84.015 85.445 ;
        RECT 84.305 85.275 84.475 85.445 ;
        RECT 84.765 85.275 84.935 85.445 ;
        RECT 85.225 85.275 85.395 85.445 ;
        RECT 85.685 85.275 85.855 85.445 ;
        RECT 86.145 85.275 86.315 85.445 ;
        RECT 86.605 85.275 86.775 85.445 ;
        RECT 87.065 85.275 87.235 85.445 ;
        RECT 87.525 85.275 87.695 85.445 ;
        RECT 87.985 85.275 88.155 85.445 ;
        RECT 88.445 85.275 88.615 85.445 ;
        RECT 88.905 85.275 89.075 85.445 ;
        RECT 89.365 85.275 89.535 85.445 ;
        RECT 89.825 85.275 89.995 85.445 ;
        RECT 90.285 85.275 90.455 85.445 ;
        RECT 90.745 85.275 90.915 85.445 ;
        RECT 91.205 85.275 91.375 85.445 ;
        RECT 91.665 85.275 91.835 85.445 ;
        RECT 92.125 85.275 92.295 85.445 ;
        RECT 92.585 85.275 92.755 85.445 ;
        RECT 93.045 85.275 93.215 85.445 ;
        RECT 93.505 85.275 93.675 85.445 ;
        RECT 93.965 85.275 94.135 85.445 ;
        RECT 94.425 85.275 94.595 85.445 ;
        RECT 94.885 85.275 95.055 85.445 ;
        RECT 95.345 85.275 95.515 85.445 ;
        RECT 95.805 85.275 95.975 85.445 ;
        RECT 96.265 85.275 96.435 85.445 ;
        RECT 96.725 85.275 96.895 85.445 ;
        RECT 97.185 85.275 97.355 85.445 ;
        RECT 97.645 85.275 97.815 85.445 ;
        RECT 98.105 85.275 98.275 85.445 ;
        RECT 98.565 85.275 98.735 85.445 ;
        RECT 99.025 85.275 99.195 85.445 ;
        RECT 99.485 85.275 99.655 85.445 ;
        RECT 99.945 85.275 100.115 85.445 ;
        RECT 100.405 85.275 100.575 85.445 ;
        RECT 100.865 85.275 101.035 85.445 ;
        RECT 101.325 85.275 101.495 85.445 ;
        RECT 101.785 85.275 101.955 85.445 ;
        RECT 102.245 85.275 102.415 85.445 ;
        RECT 102.705 85.275 102.875 85.445 ;
        RECT 103.165 85.275 103.335 85.445 ;
        RECT 103.625 85.275 103.795 85.445 ;
        RECT 104.085 85.275 104.255 85.445 ;
        RECT 104.545 85.275 104.715 85.445 ;
        RECT 105.005 85.275 105.175 85.445 ;
        RECT 105.465 85.275 105.635 85.445 ;
        RECT 105.925 85.275 106.095 85.445 ;
        RECT 106.385 85.275 106.555 85.445 ;
        RECT 106.845 85.275 107.015 85.445 ;
        RECT 107.305 85.275 107.475 85.445 ;
        RECT 107.765 85.275 107.935 85.445 ;
        RECT 108.225 85.275 108.395 85.445 ;
        RECT 108.685 85.275 108.855 85.445 ;
        RECT 109.145 85.275 109.315 85.445 ;
        RECT 109.605 85.275 109.775 85.445 ;
        RECT 110.065 85.275 110.235 85.445 ;
        RECT 110.525 85.275 110.695 85.445 ;
        RECT 110.985 85.275 111.155 85.445 ;
        RECT 111.445 85.275 111.615 85.445 ;
        RECT 111.905 85.275 112.075 85.445 ;
        RECT 112.365 85.275 112.535 85.445 ;
        RECT 112.825 85.275 112.995 85.445 ;
        RECT 113.285 85.275 113.455 85.445 ;
        RECT 113.745 85.275 113.915 85.445 ;
        RECT 114.205 85.275 114.375 85.445 ;
        RECT 114.665 85.275 114.835 85.445 ;
        RECT 115.125 85.275 115.295 85.445 ;
        RECT 115.585 85.275 115.755 85.445 ;
        RECT 116.045 85.275 116.215 85.445 ;
        RECT 116.505 85.275 116.675 85.445 ;
        RECT 116.965 85.275 117.135 85.445 ;
        RECT 117.425 85.275 117.595 85.445 ;
        RECT 117.885 85.275 118.055 85.445 ;
        RECT 118.345 85.275 118.515 85.445 ;
        RECT 118.805 85.275 118.975 85.445 ;
        RECT 119.265 85.275 119.435 85.445 ;
        RECT 119.725 85.275 119.895 85.445 ;
        RECT 120.185 85.275 120.355 85.445 ;
        RECT 120.645 85.275 120.815 85.445 ;
        RECT 121.105 85.275 121.275 85.445 ;
        RECT 121.565 85.275 121.735 85.445 ;
        RECT 122.025 85.275 122.195 85.445 ;
        RECT 122.485 85.275 122.655 85.445 ;
        RECT 122.945 85.275 123.115 85.445 ;
        RECT 123.405 85.275 123.575 85.445 ;
        RECT 123.865 85.275 124.035 85.445 ;
        RECT 124.325 85.275 124.495 85.445 ;
        RECT 124.785 85.275 124.955 85.445 ;
        RECT 125.245 85.275 125.415 85.445 ;
        RECT 125.705 85.275 125.875 85.445 ;
        RECT 126.165 85.275 126.335 85.445 ;
        RECT 126.625 85.275 126.795 85.445 ;
        RECT 127.085 85.275 127.255 85.445 ;
        RECT 127.545 85.275 127.715 85.445 ;
        RECT 128.005 85.275 128.175 85.445 ;
        RECT 128.465 85.275 128.635 85.445 ;
        RECT 128.925 85.275 129.095 85.445 ;
        RECT 129.385 85.275 129.555 85.445 ;
        RECT 129.845 85.275 130.015 85.445 ;
        RECT 130.305 85.275 130.475 85.445 ;
        RECT 130.765 85.275 130.935 85.445 ;
        RECT 131.225 85.275 131.395 85.445 ;
        RECT 131.685 85.275 131.855 85.445 ;
        RECT 132.145 85.275 132.315 85.445 ;
        RECT 132.605 85.275 132.775 85.445 ;
        RECT 133.065 85.275 133.235 85.445 ;
        RECT 133.525 85.275 133.695 85.445 ;
        RECT 133.985 85.275 134.155 85.445 ;
        RECT 45.665 79.835 45.835 80.005 ;
        RECT 46.125 79.835 46.295 80.005 ;
        RECT 46.585 79.835 46.755 80.005 ;
        RECT 47.045 79.835 47.215 80.005 ;
        RECT 47.505 79.835 47.675 80.005 ;
        RECT 47.965 79.835 48.135 80.005 ;
        RECT 48.425 79.835 48.595 80.005 ;
        RECT 48.885 79.835 49.055 80.005 ;
        RECT 49.345 79.835 49.515 80.005 ;
        RECT 49.805 79.835 49.975 80.005 ;
        RECT 50.265 79.835 50.435 80.005 ;
        RECT 50.725 79.835 50.895 80.005 ;
        RECT 51.185 79.835 51.355 80.005 ;
        RECT 51.645 79.835 51.815 80.005 ;
        RECT 52.105 79.835 52.275 80.005 ;
        RECT 52.565 79.835 52.735 80.005 ;
        RECT 53.025 79.835 53.195 80.005 ;
        RECT 53.485 79.835 53.655 80.005 ;
        RECT 53.945 79.835 54.115 80.005 ;
        RECT 54.405 79.835 54.575 80.005 ;
        RECT 54.865 79.835 55.035 80.005 ;
        RECT 55.325 79.835 55.495 80.005 ;
        RECT 55.785 79.835 55.955 80.005 ;
        RECT 56.245 79.835 56.415 80.005 ;
        RECT 56.705 79.835 56.875 80.005 ;
        RECT 57.165 79.835 57.335 80.005 ;
        RECT 57.625 79.835 57.795 80.005 ;
        RECT 58.085 79.835 58.255 80.005 ;
        RECT 58.545 79.835 58.715 80.005 ;
        RECT 59.005 79.835 59.175 80.005 ;
        RECT 59.465 79.835 59.635 80.005 ;
        RECT 59.925 79.835 60.095 80.005 ;
        RECT 60.385 79.835 60.555 80.005 ;
        RECT 60.845 79.835 61.015 80.005 ;
        RECT 61.305 79.835 61.475 80.005 ;
        RECT 61.765 79.835 61.935 80.005 ;
        RECT 62.225 79.835 62.395 80.005 ;
        RECT 62.685 79.835 62.855 80.005 ;
        RECT 63.145 79.835 63.315 80.005 ;
        RECT 63.605 79.835 63.775 80.005 ;
        RECT 64.065 79.835 64.235 80.005 ;
        RECT 64.525 79.835 64.695 80.005 ;
        RECT 64.985 79.835 65.155 80.005 ;
        RECT 65.445 79.835 65.615 80.005 ;
        RECT 65.905 79.835 66.075 80.005 ;
        RECT 66.365 79.835 66.535 80.005 ;
        RECT 66.825 79.835 66.995 80.005 ;
        RECT 67.285 79.835 67.455 80.005 ;
        RECT 67.745 79.835 67.915 80.005 ;
        RECT 68.205 79.835 68.375 80.005 ;
        RECT 68.665 79.835 68.835 80.005 ;
        RECT 69.125 79.835 69.295 80.005 ;
        RECT 69.585 79.835 69.755 80.005 ;
        RECT 70.045 79.835 70.215 80.005 ;
        RECT 70.505 79.835 70.675 80.005 ;
        RECT 70.965 79.835 71.135 80.005 ;
        RECT 71.425 79.835 71.595 80.005 ;
        RECT 71.885 79.835 72.055 80.005 ;
        RECT 72.345 79.835 72.515 80.005 ;
        RECT 72.805 79.835 72.975 80.005 ;
        RECT 73.265 79.835 73.435 80.005 ;
        RECT 73.725 79.835 73.895 80.005 ;
        RECT 74.185 79.835 74.355 80.005 ;
        RECT 74.645 79.835 74.815 80.005 ;
        RECT 75.105 79.835 75.275 80.005 ;
        RECT 75.565 79.835 75.735 80.005 ;
        RECT 76.025 79.835 76.195 80.005 ;
        RECT 76.485 79.835 76.655 80.005 ;
        RECT 76.945 79.835 77.115 80.005 ;
        RECT 77.405 79.835 77.575 80.005 ;
        RECT 77.865 79.835 78.035 80.005 ;
        RECT 78.325 79.835 78.495 80.005 ;
        RECT 78.785 79.835 78.955 80.005 ;
        RECT 79.245 79.835 79.415 80.005 ;
        RECT 79.705 79.835 79.875 80.005 ;
        RECT 80.165 79.835 80.335 80.005 ;
        RECT 80.625 79.835 80.795 80.005 ;
        RECT 81.085 79.835 81.255 80.005 ;
        RECT 81.545 79.835 81.715 80.005 ;
        RECT 82.005 79.835 82.175 80.005 ;
        RECT 82.465 79.835 82.635 80.005 ;
        RECT 82.925 79.835 83.095 80.005 ;
        RECT 83.385 79.835 83.555 80.005 ;
        RECT 83.845 79.835 84.015 80.005 ;
        RECT 84.305 79.835 84.475 80.005 ;
        RECT 84.765 79.835 84.935 80.005 ;
        RECT 85.225 79.835 85.395 80.005 ;
        RECT 85.685 79.835 85.855 80.005 ;
        RECT 86.145 79.835 86.315 80.005 ;
        RECT 86.605 79.835 86.775 80.005 ;
        RECT 87.065 79.835 87.235 80.005 ;
        RECT 87.525 79.835 87.695 80.005 ;
        RECT 87.985 79.835 88.155 80.005 ;
        RECT 88.445 79.835 88.615 80.005 ;
        RECT 88.905 79.835 89.075 80.005 ;
        RECT 89.365 79.835 89.535 80.005 ;
        RECT 89.825 79.835 89.995 80.005 ;
        RECT 90.285 79.835 90.455 80.005 ;
        RECT 90.745 79.835 90.915 80.005 ;
        RECT 91.205 79.835 91.375 80.005 ;
        RECT 91.665 79.835 91.835 80.005 ;
        RECT 92.125 79.835 92.295 80.005 ;
        RECT 92.585 79.835 92.755 80.005 ;
        RECT 93.045 79.835 93.215 80.005 ;
        RECT 93.505 79.835 93.675 80.005 ;
        RECT 93.965 79.835 94.135 80.005 ;
        RECT 94.425 79.835 94.595 80.005 ;
        RECT 94.885 79.835 95.055 80.005 ;
        RECT 95.345 79.835 95.515 80.005 ;
        RECT 95.805 79.835 95.975 80.005 ;
        RECT 96.265 79.835 96.435 80.005 ;
        RECT 96.725 79.835 96.895 80.005 ;
        RECT 97.185 79.835 97.355 80.005 ;
        RECT 97.645 79.835 97.815 80.005 ;
        RECT 98.105 79.835 98.275 80.005 ;
        RECT 98.565 79.835 98.735 80.005 ;
        RECT 99.025 79.835 99.195 80.005 ;
        RECT 99.485 79.835 99.655 80.005 ;
        RECT 99.945 79.835 100.115 80.005 ;
        RECT 100.405 79.835 100.575 80.005 ;
        RECT 100.865 79.835 101.035 80.005 ;
        RECT 101.325 79.835 101.495 80.005 ;
        RECT 101.785 79.835 101.955 80.005 ;
        RECT 102.245 79.835 102.415 80.005 ;
        RECT 102.705 79.835 102.875 80.005 ;
        RECT 103.165 79.835 103.335 80.005 ;
        RECT 103.625 79.835 103.795 80.005 ;
        RECT 104.085 79.835 104.255 80.005 ;
        RECT 104.545 79.835 104.715 80.005 ;
        RECT 105.005 79.835 105.175 80.005 ;
        RECT 105.465 79.835 105.635 80.005 ;
        RECT 105.925 79.835 106.095 80.005 ;
        RECT 106.385 79.835 106.555 80.005 ;
        RECT 106.845 79.835 107.015 80.005 ;
        RECT 107.305 79.835 107.475 80.005 ;
        RECT 107.765 79.835 107.935 80.005 ;
        RECT 108.225 79.835 108.395 80.005 ;
        RECT 108.685 79.835 108.855 80.005 ;
        RECT 109.145 79.835 109.315 80.005 ;
        RECT 109.605 79.835 109.775 80.005 ;
        RECT 110.065 79.835 110.235 80.005 ;
        RECT 110.525 79.835 110.695 80.005 ;
        RECT 110.985 79.835 111.155 80.005 ;
        RECT 111.445 79.835 111.615 80.005 ;
        RECT 111.905 79.835 112.075 80.005 ;
        RECT 112.365 79.835 112.535 80.005 ;
        RECT 112.825 79.835 112.995 80.005 ;
        RECT 113.285 79.835 113.455 80.005 ;
        RECT 113.745 79.835 113.915 80.005 ;
        RECT 114.205 79.835 114.375 80.005 ;
        RECT 114.665 79.835 114.835 80.005 ;
        RECT 115.125 79.835 115.295 80.005 ;
        RECT 115.585 79.835 115.755 80.005 ;
        RECT 116.045 79.835 116.215 80.005 ;
        RECT 116.505 79.835 116.675 80.005 ;
        RECT 116.965 79.835 117.135 80.005 ;
        RECT 117.425 79.835 117.595 80.005 ;
        RECT 117.885 79.835 118.055 80.005 ;
        RECT 118.345 79.835 118.515 80.005 ;
        RECT 118.805 79.835 118.975 80.005 ;
        RECT 119.265 79.835 119.435 80.005 ;
        RECT 119.725 79.835 119.895 80.005 ;
        RECT 120.185 79.835 120.355 80.005 ;
        RECT 120.645 79.835 120.815 80.005 ;
        RECT 121.105 79.835 121.275 80.005 ;
        RECT 121.565 79.835 121.735 80.005 ;
        RECT 122.025 79.835 122.195 80.005 ;
        RECT 122.485 79.835 122.655 80.005 ;
        RECT 122.945 79.835 123.115 80.005 ;
        RECT 123.405 79.835 123.575 80.005 ;
        RECT 123.865 79.835 124.035 80.005 ;
        RECT 124.325 79.835 124.495 80.005 ;
        RECT 124.785 79.835 124.955 80.005 ;
        RECT 125.245 79.835 125.415 80.005 ;
        RECT 125.705 79.835 125.875 80.005 ;
        RECT 126.165 79.835 126.335 80.005 ;
        RECT 126.625 79.835 126.795 80.005 ;
        RECT 127.085 79.835 127.255 80.005 ;
        RECT 127.545 79.835 127.715 80.005 ;
        RECT 128.005 79.835 128.175 80.005 ;
        RECT 128.465 79.835 128.635 80.005 ;
        RECT 128.925 79.835 129.095 80.005 ;
        RECT 129.385 79.835 129.555 80.005 ;
        RECT 129.845 79.835 130.015 80.005 ;
        RECT 130.305 79.835 130.475 80.005 ;
        RECT 130.765 79.835 130.935 80.005 ;
        RECT 131.225 79.835 131.395 80.005 ;
        RECT 131.685 79.835 131.855 80.005 ;
        RECT 132.145 79.835 132.315 80.005 ;
        RECT 132.605 79.835 132.775 80.005 ;
        RECT 133.065 79.835 133.235 80.005 ;
        RECT 133.525 79.835 133.695 80.005 ;
        RECT 133.985 79.835 134.155 80.005 ;
        RECT 45.665 74.395 45.835 74.565 ;
        RECT 46.125 74.395 46.295 74.565 ;
        RECT 46.585 74.395 46.755 74.565 ;
        RECT 47.045 74.395 47.215 74.565 ;
        RECT 47.505 74.395 47.675 74.565 ;
        RECT 47.965 74.395 48.135 74.565 ;
        RECT 48.425 74.395 48.595 74.565 ;
        RECT 48.885 74.395 49.055 74.565 ;
        RECT 49.345 74.395 49.515 74.565 ;
        RECT 49.805 74.395 49.975 74.565 ;
        RECT 50.265 74.395 50.435 74.565 ;
        RECT 50.725 74.395 50.895 74.565 ;
        RECT 51.185 74.395 51.355 74.565 ;
        RECT 51.645 74.395 51.815 74.565 ;
        RECT 52.105 74.395 52.275 74.565 ;
        RECT 52.565 74.395 52.735 74.565 ;
        RECT 53.025 74.395 53.195 74.565 ;
        RECT 53.485 74.395 53.655 74.565 ;
        RECT 53.945 74.395 54.115 74.565 ;
        RECT 54.405 74.395 54.575 74.565 ;
        RECT 54.865 74.395 55.035 74.565 ;
        RECT 55.325 74.395 55.495 74.565 ;
        RECT 55.785 74.395 55.955 74.565 ;
        RECT 56.245 74.395 56.415 74.565 ;
        RECT 56.705 74.395 56.875 74.565 ;
        RECT 57.165 74.395 57.335 74.565 ;
        RECT 57.625 74.395 57.795 74.565 ;
        RECT 58.085 74.395 58.255 74.565 ;
        RECT 58.545 74.395 58.715 74.565 ;
        RECT 59.005 74.395 59.175 74.565 ;
        RECT 59.465 74.395 59.635 74.565 ;
        RECT 59.925 74.395 60.095 74.565 ;
        RECT 60.385 74.395 60.555 74.565 ;
        RECT 60.845 74.395 61.015 74.565 ;
        RECT 61.305 74.395 61.475 74.565 ;
        RECT 61.765 74.395 61.935 74.565 ;
        RECT 62.225 74.395 62.395 74.565 ;
        RECT 62.685 74.395 62.855 74.565 ;
        RECT 63.145 74.395 63.315 74.565 ;
        RECT 63.605 74.395 63.775 74.565 ;
        RECT 64.065 74.395 64.235 74.565 ;
        RECT 64.525 74.395 64.695 74.565 ;
        RECT 64.985 74.395 65.155 74.565 ;
        RECT 65.445 74.395 65.615 74.565 ;
        RECT 65.905 74.395 66.075 74.565 ;
        RECT 66.365 74.395 66.535 74.565 ;
        RECT 66.825 74.395 66.995 74.565 ;
        RECT 67.285 74.395 67.455 74.565 ;
        RECT 67.745 74.395 67.915 74.565 ;
        RECT 68.205 74.395 68.375 74.565 ;
        RECT 68.665 74.395 68.835 74.565 ;
        RECT 69.125 74.395 69.295 74.565 ;
        RECT 69.585 74.395 69.755 74.565 ;
        RECT 70.045 74.395 70.215 74.565 ;
        RECT 70.505 74.395 70.675 74.565 ;
        RECT 70.965 74.395 71.135 74.565 ;
        RECT 71.425 74.395 71.595 74.565 ;
        RECT 71.885 74.395 72.055 74.565 ;
        RECT 72.345 74.395 72.515 74.565 ;
        RECT 72.805 74.395 72.975 74.565 ;
        RECT 73.265 74.395 73.435 74.565 ;
        RECT 73.725 74.395 73.895 74.565 ;
        RECT 74.185 74.395 74.355 74.565 ;
        RECT 74.645 74.395 74.815 74.565 ;
        RECT 75.105 74.395 75.275 74.565 ;
        RECT 75.565 74.395 75.735 74.565 ;
        RECT 76.025 74.395 76.195 74.565 ;
        RECT 76.485 74.395 76.655 74.565 ;
        RECT 76.945 74.395 77.115 74.565 ;
        RECT 77.405 74.395 77.575 74.565 ;
        RECT 77.865 74.395 78.035 74.565 ;
        RECT 78.325 74.395 78.495 74.565 ;
        RECT 78.785 74.395 78.955 74.565 ;
        RECT 79.245 74.395 79.415 74.565 ;
        RECT 79.705 74.395 79.875 74.565 ;
        RECT 80.165 74.395 80.335 74.565 ;
        RECT 80.625 74.395 80.795 74.565 ;
        RECT 81.085 74.395 81.255 74.565 ;
        RECT 81.545 74.395 81.715 74.565 ;
        RECT 82.005 74.395 82.175 74.565 ;
        RECT 82.465 74.395 82.635 74.565 ;
        RECT 82.925 74.395 83.095 74.565 ;
        RECT 83.385 74.395 83.555 74.565 ;
        RECT 83.845 74.395 84.015 74.565 ;
        RECT 84.305 74.395 84.475 74.565 ;
        RECT 84.765 74.395 84.935 74.565 ;
        RECT 85.225 74.395 85.395 74.565 ;
        RECT 85.685 74.395 85.855 74.565 ;
        RECT 86.145 74.395 86.315 74.565 ;
        RECT 86.605 74.395 86.775 74.565 ;
        RECT 87.065 74.395 87.235 74.565 ;
        RECT 87.525 74.395 87.695 74.565 ;
        RECT 87.985 74.395 88.155 74.565 ;
        RECT 88.445 74.395 88.615 74.565 ;
        RECT 88.905 74.395 89.075 74.565 ;
        RECT 89.365 74.395 89.535 74.565 ;
        RECT 89.825 74.395 89.995 74.565 ;
        RECT 90.285 74.395 90.455 74.565 ;
        RECT 90.745 74.395 90.915 74.565 ;
        RECT 91.205 74.395 91.375 74.565 ;
        RECT 91.665 74.395 91.835 74.565 ;
        RECT 92.125 74.395 92.295 74.565 ;
        RECT 92.585 74.395 92.755 74.565 ;
        RECT 93.045 74.395 93.215 74.565 ;
        RECT 93.505 74.395 93.675 74.565 ;
        RECT 93.965 74.395 94.135 74.565 ;
        RECT 94.425 74.395 94.595 74.565 ;
        RECT 94.885 74.395 95.055 74.565 ;
        RECT 95.345 74.395 95.515 74.565 ;
        RECT 95.805 74.395 95.975 74.565 ;
        RECT 96.265 74.395 96.435 74.565 ;
        RECT 96.725 74.395 96.895 74.565 ;
        RECT 97.185 74.395 97.355 74.565 ;
        RECT 97.645 74.395 97.815 74.565 ;
        RECT 98.105 74.395 98.275 74.565 ;
        RECT 98.565 74.395 98.735 74.565 ;
        RECT 99.025 74.395 99.195 74.565 ;
        RECT 99.485 74.395 99.655 74.565 ;
        RECT 99.945 74.395 100.115 74.565 ;
        RECT 100.405 74.395 100.575 74.565 ;
        RECT 100.865 74.395 101.035 74.565 ;
        RECT 101.325 74.395 101.495 74.565 ;
        RECT 101.785 74.395 101.955 74.565 ;
        RECT 102.245 74.395 102.415 74.565 ;
        RECT 102.705 74.395 102.875 74.565 ;
        RECT 103.165 74.395 103.335 74.565 ;
        RECT 103.625 74.395 103.795 74.565 ;
        RECT 104.085 74.395 104.255 74.565 ;
        RECT 104.545 74.395 104.715 74.565 ;
        RECT 105.005 74.395 105.175 74.565 ;
        RECT 105.465 74.395 105.635 74.565 ;
        RECT 105.925 74.395 106.095 74.565 ;
        RECT 106.385 74.395 106.555 74.565 ;
        RECT 106.845 74.395 107.015 74.565 ;
        RECT 107.305 74.395 107.475 74.565 ;
        RECT 107.765 74.395 107.935 74.565 ;
        RECT 108.225 74.395 108.395 74.565 ;
        RECT 108.685 74.395 108.855 74.565 ;
        RECT 109.145 74.395 109.315 74.565 ;
        RECT 109.605 74.395 109.775 74.565 ;
        RECT 110.065 74.395 110.235 74.565 ;
        RECT 110.525 74.395 110.695 74.565 ;
        RECT 110.985 74.395 111.155 74.565 ;
        RECT 111.445 74.395 111.615 74.565 ;
        RECT 111.905 74.395 112.075 74.565 ;
        RECT 112.365 74.395 112.535 74.565 ;
        RECT 112.825 74.395 112.995 74.565 ;
        RECT 113.285 74.395 113.455 74.565 ;
        RECT 113.745 74.395 113.915 74.565 ;
        RECT 114.205 74.395 114.375 74.565 ;
        RECT 114.665 74.395 114.835 74.565 ;
        RECT 115.125 74.395 115.295 74.565 ;
        RECT 115.585 74.395 115.755 74.565 ;
        RECT 116.045 74.395 116.215 74.565 ;
        RECT 116.505 74.395 116.675 74.565 ;
        RECT 116.965 74.395 117.135 74.565 ;
        RECT 117.425 74.395 117.595 74.565 ;
        RECT 117.885 74.395 118.055 74.565 ;
        RECT 118.345 74.395 118.515 74.565 ;
        RECT 118.805 74.395 118.975 74.565 ;
        RECT 119.265 74.395 119.435 74.565 ;
        RECT 119.725 74.395 119.895 74.565 ;
        RECT 120.185 74.395 120.355 74.565 ;
        RECT 120.645 74.395 120.815 74.565 ;
        RECT 121.105 74.395 121.275 74.565 ;
        RECT 121.565 74.395 121.735 74.565 ;
        RECT 122.025 74.395 122.195 74.565 ;
        RECT 122.485 74.395 122.655 74.565 ;
        RECT 122.945 74.395 123.115 74.565 ;
        RECT 123.405 74.395 123.575 74.565 ;
        RECT 123.865 74.395 124.035 74.565 ;
        RECT 124.325 74.395 124.495 74.565 ;
        RECT 124.785 74.395 124.955 74.565 ;
        RECT 125.245 74.395 125.415 74.565 ;
        RECT 125.705 74.395 125.875 74.565 ;
        RECT 126.165 74.395 126.335 74.565 ;
        RECT 126.625 74.395 126.795 74.565 ;
        RECT 127.085 74.395 127.255 74.565 ;
        RECT 127.545 74.395 127.715 74.565 ;
        RECT 128.005 74.395 128.175 74.565 ;
        RECT 128.465 74.395 128.635 74.565 ;
        RECT 128.925 74.395 129.095 74.565 ;
        RECT 129.385 74.395 129.555 74.565 ;
        RECT 129.845 74.395 130.015 74.565 ;
        RECT 130.305 74.395 130.475 74.565 ;
        RECT 130.765 74.395 130.935 74.565 ;
        RECT 131.225 74.395 131.395 74.565 ;
        RECT 131.685 74.395 131.855 74.565 ;
        RECT 132.145 74.395 132.315 74.565 ;
        RECT 132.605 74.395 132.775 74.565 ;
        RECT 133.065 74.395 133.235 74.565 ;
        RECT 133.525 74.395 133.695 74.565 ;
        RECT 133.985 74.395 134.155 74.565 ;
        RECT 45.665 68.955 45.835 69.125 ;
        RECT 46.125 68.955 46.295 69.125 ;
        RECT 46.585 68.955 46.755 69.125 ;
        RECT 47.045 68.955 47.215 69.125 ;
        RECT 47.505 68.955 47.675 69.125 ;
        RECT 47.965 68.955 48.135 69.125 ;
        RECT 48.425 68.955 48.595 69.125 ;
        RECT 48.885 68.955 49.055 69.125 ;
        RECT 49.345 68.955 49.515 69.125 ;
        RECT 49.805 68.955 49.975 69.125 ;
        RECT 50.265 68.955 50.435 69.125 ;
        RECT 50.725 68.955 50.895 69.125 ;
        RECT 51.185 68.955 51.355 69.125 ;
        RECT 51.645 68.955 51.815 69.125 ;
        RECT 52.105 68.955 52.275 69.125 ;
        RECT 52.565 68.955 52.735 69.125 ;
        RECT 53.025 68.955 53.195 69.125 ;
        RECT 53.485 68.955 53.655 69.125 ;
        RECT 53.945 68.955 54.115 69.125 ;
        RECT 54.405 68.955 54.575 69.125 ;
        RECT 54.865 68.955 55.035 69.125 ;
        RECT 55.325 68.955 55.495 69.125 ;
        RECT 55.785 68.955 55.955 69.125 ;
        RECT 56.245 68.955 56.415 69.125 ;
        RECT 56.705 68.955 56.875 69.125 ;
        RECT 57.165 68.955 57.335 69.125 ;
        RECT 57.625 68.955 57.795 69.125 ;
        RECT 58.085 68.955 58.255 69.125 ;
        RECT 58.545 68.955 58.715 69.125 ;
        RECT 59.005 68.955 59.175 69.125 ;
        RECT 59.465 68.955 59.635 69.125 ;
        RECT 59.925 68.955 60.095 69.125 ;
        RECT 60.385 68.955 60.555 69.125 ;
        RECT 60.845 68.955 61.015 69.125 ;
        RECT 61.305 68.955 61.475 69.125 ;
        RECT 61.765 68.955 61.935 69.125 ;
        RECT 62.225 68.955 62.395 69.125 ;
        RECT 62.685 68.955 62.855 69.125 ;
        RECT 63.145 68.955 63.315 69.125 ;
        RECT 63.605 68.955 63.775 69.125 ;
        RECT 64.065 68.955 64.235 69.125 ;
        RECT 64.525 68.955 64.695 69.125 ;
        RECT 64.985 68.955 65.155 69.125 ;
        RECT 65.445 68.955 65.615 69.125 ;
        RECT 65.905 68.955 66.075 69.125 ;
        RECT 66.365 68.955 66.535 69.125 ;
        RECT 66.825 68.955 66.995 69.125 ;
        RECT 67.285 68.955 67.455 69.125 ;
        RECT 67.745 68.955 67.915 69.125 ;
        RECT 68.205 68.955 68.375 69.125 ;
        RECT 68.665 68.955 68.835 69.125 ;
        RECT 69.125 68.955 69.295 69.125 ;
        RECT 69.585 68.955 69.755 69.125 ;
        RECT 70.045 68.955 70.215 69.125 ;
        RECT 70.505 68.955 70.675 69.125 ;
        RECT 70.965 68.955 71.135 69.125 ;
        RECT 71.425 68.955 71.595 69.125 ;
        RECT 71.885 68.955 72.055 69.125 ;
        RECT 72.345 68.955 72.515 69.125 ;
        RECT 72.805 68.955 72.975 69.125 ;
        RECT 73.265 68.955 73.435 69.125 ;
        RECT 73.725 68.955 73.895 69.125 ;
        RECT 74.185 68.955 74.355 69.125 ;
        RECT 74.645 68.955 74.815 69.125 ;
        RECT 75.105 68.955 75.275 69.125 ;
        RECT 75.565 68.955 75.735 69.125 ;
        RECT 76.025 68.955 76.195 69.125 ;
        RECT 76.485 68.955 76.655 69.125 ;
        RECT 76.945 68.955 77.115 69.125 ;
        RECT 77.405 68.955 77.575 69.125 ;
        RECT 77.865 68.955 78.035 69.125 ;
        RECT 78.325 68.955 78.495 69.125 ;
        RECT 78.785 68.955 78.955 69.125 ;
        RECT 79.245 68.955 79.415 69.125 ;
        RECT 79.705 68.955 79.875 69.125 ;
        RECT 80.165 68.955 80.335 69.125 ;
        RECT 80.625 68.955 80.795 69.125 ;
        RECT 81.085 68.955 81.255 69.125 ;
        RECT 81.545 68.955 81.715 69.125 ;
        RECT 82.005 68.955 82.175 69.125 ;
        RECT 82.465 68.955 82.635 69.125 ;
        RECT 82.925 68.955 83.095 69.125 ;
        RECT 83.385 68.955 83.555 69.125 ;
        RECT 83.845 68.955 84.015 69.125 ;
        RECT 84.305 68.955 84.475 69.125 ;
        RECT 84.765 68.955 84.935 69.125 ;
        RECT 85.225 68.955 85.395 69.125 ;
        RECT 85.685 68.955 85.855 69.125 ;
        RECT 86.145 68.955 86.315 69.125 ;
        RECT 86.605 68.955 86.775 69.125 ;
        RECT 87.065 68.955 87.235 69.125 ;
        RECT 87.525 68.955 87.695 69.125 ;
        RECT 87.985 68.955 88.155 69.125 ;
        RECT 88.445 68.955 88.615 69.125 ;
        RECT 88.905 68.955 89.075 69.125 ;
        RECT 89.365 68.955 89.535 69.125 ;
        RECT 89.825 68.955 89.995 69.125 ;
        RECT 90.285 68.955 90.455 69.125 ;
        RECT 90.745 68.955 90.915 69.125 ;
        RECT 91.205 68.955 91.375 69.125 ;
        RECT 91.665 68.955 91.835 69.125 ;
        RECT 92.125 68.955 92.295 69.125 ;
        RECT 92.585 68.955 92.755 69.125 ;
        RECT 93.045 68.955 93.215 69.125 ;
        RECT 93.505 68.955 93.675 69.125 ;
        RECT 93.965 68.955 94.135 69.125 ;
        RECT 94.425 68.955 94.595 69.125 ;
        RECT 94.885 68.955 95.055 69.125 ;
        RECT 95.345 68.955 95.515 69.125 ;
        RECT 95.805 68.955 95.975 69.125 ;
        RECT 96.265 68.955 96.435 69.125 ;
        RECT 96.725 68.955 96.895 69.125 ;
        RECT 97.185 68.955 97.355 69.125 ;
        RECT 97.645 68.955 97.815 69.125 ;
        RECT 98.105 68.955 98.275 69.125 ;
        RECT 98.565 68.955 98.735 69.125 ;
        RECT 99.025 68.955 99.195 69.125 ;
        RECT 99.485 68.955 99.655 69.125 ;
        RECT 99.945 68.955 100.115 69.125 ;
        RECT 100.405 68.955 100.575 69.125 ;
        RECT 100.865 68.955 101.035 69.125 ;
        RECT 101.325 68.955 101.495 69.125 ;
        RECT 101.785 68.955 101.955 69.125 ;
        RECT 102.245 68.955 102.415 69.125 ;
        RECT 102.705 68.955 102.875 69.125 ;
        RECT 103.165 68.955 103.335 69.125 ;
        RECT 103.625 68.955 103.795 69.125 ;
        RECT 104.085 68.955 104.255 69.125 ;
        RECT 104.545 68.955 104.715 69.125 ;
        RECT 105.005 68.955 105.175 69.125 ;
        RECT 105.465 68.955 105.635 69.125 ;
        RECT 105.925 68.955 106.095 69.125 ;
        RECT 106.385 68.955 106.555 69.125 ;
        RECT 106.845 68.955 107.015 69.125 ;
        RECT 107.305 68.955 107.475 69.125 ;
        RECT 107.765 68.955 107.935 69.125 ;
        RECT 108.225 68.955 108.395 69.125 ;
        RECT 108.685 68.955 108.855 69.125 ;
        RECT 109.145 68.955 109.315 69.125 ;
        RECT 109.605 68.955 109.775 69.125 ;
        RECT 110.065 68.955 110.235 69.125 ;
        RECT 110.525 68.955 110.695 69.125 ;
        RECT 110.985 68.955 111.155 69.125 ;
        RECT 111.445 68.955 111.615 69.125 ;
        RECT 111.905 68.955 112.075 69.125 ;
        RECT 112.365 68.955 112.535 69.125 ;
        RECT 112.825 68.955 112.995 69.125 ;
        RECT 113.285 68.955 113.455 69.125 ;
        RECT 113.745 68.955 113.915 69.125 ;
        RECT 114.205 68.955 114.375 69.125 ;
        RECT 114.665 68.955 114.835 69.125 ;
        RECT 115.125 68.955 115.295 69.125 ;
        RECT 115.585 68.955 115.755 69.125 ;
        RECT 116.045 68.955 116.215 69.125 ;
        RECT 116.505 68.955 116.675 69.125 ;
        RECT 116.965 68.955 117.135 69.125 ;
        RECT 117.425 68.955 117.595 69.125 ;
        RECT 117.885 68.955 118.055 69.125 ;
        RECT 118.345 68.955 118.515 69.125 ;
        RECT 118.805 68.955 118.975 69.125 ;
        RECT 119.265 68.955 119.435 69.125 ;
        RECT 119.725 68.955 119.895 69.125 ;
        RECT 120.185 68.955 120.355 69.125 ;
        RECT 120.645 68.955 120.815 69.125 ;
        RECT 121.105 68.955 121.275 69.125 ;
        RECT 121.565 68.955 121.735 69.125 ;
        RECT 122.025 68.955 122.195 69.125 ;
        RECT 122.485 68.955 122.655 69.125 ;
        RECT 122.945 68.955 123.115 69.125 ;
        RECT 123.405 68.955 123.575 69.125 ;
        RECT 123.865 68.955 124.035 69.125 ;
        RECT 124.325 68.955 124.495 69.125 ;
        RECT 124.785 68.955 124.955 69.125 ;
        RECT 125.245 68.955 125.415 69.125 ;
        RECT 125.705 68.955 125.875 69.125 ;
        RECT 126.165 68.955 126.335 69.125 ;
        RECT 126.625 68.955 126.795 69.125 ;
        RECT 127.085 68.955 127.255 69.125 ;
        RECT 127.545 68.955 127.715 69.125 ;
        RECT 128.005 68.955 128.175 69.125 ;
        RECT 128.465 68.955 128.635 69.125 ;
        RECT 128.925 68.955 129.095 69.125 ;
        RECT 129.385 68.955 129.555 69.125 ;
        RECT 129.845 68.955 130.015 69.125 ;
        RECT 130.305 68.955 130.475 69.125 ;
        RECT 130.765 68.955 130.935 69.125 ;
        RECT 131.225 68.955 131.395 69.125 ;
        RECT 131.685 68.955 131.855 69.125 ;
        RECT 132.145 68.955 132.315 69.125 ;
        RECT 132.605 68.955 132.775 69.125 ;
        RECT 133.065 68.955 133.235 69.125 ;
        RECT 133.525 68.955 133.695 69.125 ;
        RECT 133.985 68.955 134.155 69.125 ;
        RECT 45.665 63.515 45.835 63.685 ;
        RECT 46.125 63.515 46.295 63.685 ;
        RECT 46.585 63.515 46.755 63.685 ;
        RECT 47.045 63.515 47.215 63.685 ;
        RECT 47.505 63.515 47.675 63.685 ;
        RECT 47.965 63.515 48.135 63.685 ;
        RECT 48.425 63.515 48.595 63.685 ;
        RECT 48.885 63.515 49.055 63.685 ;
        RECT 49.345 63.515 49.515 63.685 ;
        RECT 49.805 63.515 49.975 63.685 ;
        RECT 50.265 63.515 50.435 63.685 ;
        RECT 50.725 63.515 50.895 63.685 ;
        RECT 51.185 63.515 51.355 63.685 ;
        RECT 51.645 63.515 51.815 63.685 ;
        RECT 52.105 63.515 52.275 63.685 ;
        RECT 52.565 63.515 52.735 63.685 ;
        RECT 53.025 63.515 53.195 63.685 ;
        RECT 53.485 63.515 53.655 63.685 ;
        RECT 53.945 63.515 54.115 63.685 ;
        RECT 54.405 63.515 54.575 63.685 ;
        RECT 54.865 63.515 55.035 63.685 ;
        RECT 55.325 63.515 55.495 63.685 ;
        RECT 55.785 63.515 55.955 63.685 ;
        RECT 56.245 63.515 56.415 63.685 ;
        RECT 56.705 63.515 56.875 63.685 ;
        RECT 57.165 63.515 57.335 63.685 ;
        RECT 57.625 63.515 57.795 63.685 ;
        RECT 58.085 63.515 58.255 63.685 ;
        RECT 58.545 63.515 58.715 63.685 ;
        RECT 59.005 63.515 59.175 63.685 ;
        RECT 59.465 63.515 59.635 63.685 ;
        RECT 59.925 63.515 60.095 63.685 ;
        RECT 60.385 63.515 60.555 63.685 ;
        RECT 60.845 63.515 61.015 63.685 ;
        RECT 61.305 63.515 61.475 63.685 ;
        RECT 61.765 63.515 61.935 63.685 ;
        RECT 62.225 63.515 62.395 63.685 ;
        RECT 62.685 63.515 62.855 63.685 ;
        RECT 63.145 63.515 63.315 63.685 ;
        RECT 63.605 63.515 63.775 63.685 ;
        RECT 64.065 63.515 64.235 63.685 ;
        RECT 64.525 63.515 64.695 63.685 ;
        RECT 64.985 63.515 65.155 63.685 ;
        RECT 65.445 63.515 65.615 63.685 ;
        RECT 65.905 63.515 66.075 63.685 ;
        RECT 66.365 63.515 66.535 63.685 ;
        RECT 66.825 63.515 66.995 63.685 ;
        RECT 67.285 63.515 67.455 63.685 ;
        RECT 67.745 63.515 67.915 63.685 ;
        RECT 68.205 63.515 68.375 63.685 ;
        RECT 68.665 63.515 68.835 63.685 ;
        RECT 69.125 63.515 69.295 63.685 ;
        RECT 69.585 63.515 69.755 63.685 ;
        RECT 70.045 63.515 70.215 63.685 ;
        RECT 70.505 63.515 70.675 63.685 ;
        RECT 70.965 63.515 71.135 63.685 ;
        RECT 71.425 63.515 71.595 63.685 ;
        RECT 71.885 63.515 72.055 63.685 ;
        RECT 72.345 63.515 72.515 63.685 ;
        RECT 72.805 63.515 72.975 63.685 ;
        RECT 73.265 63.515 73.435 63.685 ;
        RECT 73.725 63.515 73.895 63.685 ;
        RECT 74.185 63.515 74.355 63.685 ;
        RECT 74.645 63.515 74.815 63.685 ;
        RECT 75.105 63.515 75.275 63.685 ;
        RECT 75.565 63.515 75.735 63.685 ;
        RECT 76.025 63.515 76.195 63.685 ;
        RECT 76.485 63.515 76.655 63.685 ;
        RECT 76.945 63.515 77.115 63.685 ;
        RECT 77.405 63.515 77.575 63.685 ;
        RECT 77.865 63.515 78.035 63.685 ;
        RECT 78.325 63.515 78.495 63.685 ;
        RECT 78.785 63.515 78.955 63.685 ;
        RECT 79.245 63.515 79.415 63.685 ;
        RECT 79.705 63.515 79.875 63.685 ;
        RECT 80.165 63.515 80.335 63.685 ;
        RECT 80.625 63.515 80.795 63.685 ;
        RECT 81.085 63.515 81.255 63.685 ;
        RECT 81.545 63.515 81.715 63.685 ;
        RECT 82.005 63.515 82.175 63.685 ;
        RECT 82.465 63.515 82.635 63.685 ;
        RECT 82.925 63.515 83.095 63.685 ;
        RECT 83.385 63.515 83.555 63.685 ;
        RECT 83.845 63.515 84.015 63.685 ;
        RECT 84.305 63.515 84.475 63.685 ;
        RECT 84.765 63.515 84.935 63.685 ;
        RECT 85.225 63.515 85.395 63.685 ;
        RECT 85.685 63.515 85.855 63.685 ;
        RECT 86.145 63.515 86.315 63.685 ;
        RECT 86.605 63.515 86.775 63.685 ;
        RECT 87.065 63.515 87.235 63.685 ;
        RECT 87.525 63.515 87.695 63.685 ;
        RECT 87.985 63.515 88.155 63.685 ;
        RECT 88.445 63.515 88.615 63.685 ;
        RECT 88.905 63.515 89.075 63.685 ;
        RECT 89.365 63.515 89.535 63.685 ;
        RECT 89.825 63.515 89.995 63.685 ;
        RECT 90.285 63.515 90.455 63.685 ;
        RECT 90.745 63.515 90.915 63.685 ;
        RECT 91.205 63.515 91.375 63.685 ;
        RECT 91.665 63.515 91.835 63.685 ;
        RECT 92.125 63.515 92.295 63.685 ;
        RECT 92.585 63.515 92.755 63.685 ;
        RECT 93.045 63.515 93.215 63.685 ;
        RECT 93.505 63.515 93.675 63.685 ;
        RECT 93.965 63.515 94.135 63.685 ;
        RECT 94.425 63.515 94.595 63.685 ;
        RECT 94.885 63.515 95.055 63.685 ;
        RECT 95.345 63.515 95.515 63.685 ;
        RECT 95.805 63.515 95.975 63.685 ;
        RECT 96.265 63.515 96.435 63.685 ;
        RECT 96.725 63.515 96.895 63.685 ;
        RECT 97.185 63.515 97.355 63.685 ;
        RECT 97.645 63.515 97.815 63.685 ;
        RECT 98.105 63.515 98.275 63.685 ;
        RECT 98.565 63.515 98.735 63.685 ;
        RECT 99.025 63.515 99.195 63.685 ;
        RECT 99.485 63.515 99.655 63.685 ;
        RECT 99.945 63.515 100.115 63.685 ;
        RECT 100.405 63.515 100.575 63.685 ;
        RECT 100.865 63.515 101.035 63.685 ;
        RECT 101.325 63.515 101.495 63.685 ;
        RECT 101.785 63.515 101.955 63.685 ;
        RECT 102.245 63.515 102.415 63.685 ;
        RECT 102.705 63.515 102.875 63.685 ;
        RECT 103.165 63.515 103.335 63.685 ;
        RECT 103.625 63.515 103.795 63.685 ;
        RECT 104.085 63.515 104.255 63.685 ;
        RECT 104.545 63.515 104.715 63.685 ;
        RECT 105.005 63.515 105.175 63.685 ;
        RECT 105.465 63.515 105.635 63.685 ;
        RECT 105.925 63.515 106.095 63.685 ;
        RECT 106.385 63.515 106.555 63.685 ;
        RECT 106.845 63.515 107.015 63.685 ;
        RECT 107.305 63.515 107.475 63.685 ;
        RECT 107.765 63.515 107.935 63.685 ;
        RECT 108.225 63.515 108.395 63.685 ;
        RECT 108.685 63.515 108.855 63.685 ;
        RECT 109.145 63.515 109.315 63.685 ;
        RECT 109.605 63.515 109.775 63.685 ;
        RECT 110.065 63.515 110.235 63.685 ;
        RECT 110.525 63.515 110.695 63.685 ;
        RECT 110.985 63.515 111.155 63.685 ;
        RECT 111.445 63.515 111.615 63.685 ;
        RECT 111.905 63.515 112.075 63.685 ;
        RECT 112.365 63.515 112.535 63.685 ;
        RECT 112.825 63.515 112.995 63.685 ;
        RECT 113.285 63.515 113.455 63.685 ;
        RECT 113.745 63.515 113.915 63.685 ;
        RECT 114.205 63.515 114.375 63.685 ;
        RECT 114.665 63.515 114.835 63.685 ;
        RECT 115.125 63.515 115.295 63.685 ;
        RECT 115.585 63.515 115.755 63.685 ;
        RECT 116.045 63.515 116.215 63.685 ;
        RECT 116.505 63.515 116.675 63.685 ;
        RECT 116.965 63.515 117.135 63.685 ;
        RECT 117.425 63.515 117.595 63.685 ;
        RECT 117.885 63.515 118.055 63.685 ;
        RECT 118.345 63.515 118.515 63.685 ;
        RECT 118.805 63.515 118.975 63.685 ;
        RECT 119.265 63.515 119.435 63.685 ;
        RECT 119.725 63.515 119.895 63.685 ;
        RECT 120.185 63.515 120.355 63.685 ;
        RECT 120.645 63.515 120.815 63.685 ;
        RECT 121.105 63.515 121.275 63.685 ;
        RECT 121.565 63.515 121.735 63.685 ;
        RECT 122.025 63.515 122.195 63.685 ;
        RECT 122.485 63.515 122.655 63.685 ;
        RECT 122.945 63.515 123.115 63.685 ;
        RECT 123.405 63.515 123.575 63.685 ;
        RECT 123.865 63.515 124.035 63.685 ;
        RECT 124.325 63.515 124.495 63.685 ;
        RECT 124.785 63.515 124.955 63.685 ;
        RECT 125.245 63.515 125.415 63.685 ;
        RECT 125.705 63.515 125.875 63.685 ;
        RECT 126.165 63.515 126.335 63.685 ;
        RECT 126.625 63.515 126.795 63.685 ;
        RECT 127.085 63.515 127.255 63.685 ;
        RECT 127.545 63.515 127.715 63.685 ;
        RECT 128.005 63.515 128.175 63.685 ;
        RECT 128.465 63.515 128.635 63.685 ;
        RECT 128.925 63.515 129.095 63.685 ;
        RECT 129.385 63.515 129.555 63.685 ;
        RECT 129.845 63.515 130.015 63.685 ;
        RECT 130.305 63.515 130.475 63.685 ;
        RECT 130.765 63.515 130.935 63.685 ;
        RECT 131.225 63.515 131.395 63.685 ;
        RECT 131.685 63.515 131.855 63.685 ;
        RECT 132.145 63.515 132.315 63.685 ;
        RECT 132.605 63.515 132.775 63.685 ;
        RECT 133.065 63.515 133.235 63.685 ;
        RECT 133.525 63.515 133.695 63.685 ;
        RECT 133.985 63.515 134.155 63.685 ;
      LAYER met1 ;
        RECT 45.520 134.080 134.300 134.560 ;
        RECT 45.520 128.640 134.300 129.120 ;
        RECT 45.520 123.200 134.300 123.680 ;
        RECT 45.520 117.760 134.300 118.240 ;
        RECT 45.520 112.320 134.300 112.800 ;
        RECT 45.520 106.880 134.300 107.360 ;
        RECT 45.520 101.440 134.300 101.920 ;
        RECT 45.520 96.000 134.300 96.480 ;
        RECT 45.520 90.560 134.300 91.040 ;
        RECT 45.520 85.120 134.300 85.600 ;
        RECT 45.520 79.680 134.300 80.160 ;
        RECT 45.520 74.240 134.300 74.720 ;
        RECT 45.520 68.800 134.300 69.280 ;
        RECT 45.520 63.360 134.300 63.840 ;
      LAYER via ;
        RECT 55.845 134.190 56.105 134.450 ;
        RECT 56.165 134.190 56.425 134.450 ;
        RECT 56.485 134.190 56.745 134.450 ;
        RECT 56.805 134.190 57.065 134.450 ;
        RECT 57.125 134.190 57.385 134.450 ;
        RECT 78.040 134.190 78.300 134.450 ;
        RECT 78.360 134.190 78.620 134.450 ;
        RECT 78.680 134.190 78.940 134.450 ;
        RECT 79.000 134.190 79.260 134.450 ;
        RECT 79.320 134.190 79.580 134.450 ;
        RECT 100.235 134.190 100.495 134.450 ;
        RECT 100.555 134.190 100.815 134.450 ;
        RECT 100.875 134.190 101.135 134.450 ;
        RECT 101.195 134.190 101.455 134.450 ;
        RECT 101.515 134.190 101.775 134.450 ;
        RECT 122.430 134.190 122.690 134.450 ;
        RECT 122.750 134.190 123.010 134.450 ;
        RECT 123.070 134.190 123.330 134.450 ;
        RECT 123.390 134.190 123.650 134.450 ;
        RECT 123.710 134.190 123.970 134.450 ;
        RECT 55.845 128.750 56.105 129.010 ;
        RECT 56.165 128.750 56.425 129.010 ;
        RECT 56.485 128.750 56.745 129.010 ;
        RECT 56.805 128.750 57.065 129.010 ;
        RECT 57.125 128.750 57.385 129.010 ;
        RECT 78.040 128.750 78.300 129.010 ;
        RECT 78.360 128.750 78.620 129.010 ;
        RECT 78.680 128.750 78.940 129.010 ;
        RECT 79.000 128.750 79.260 129.010 ;
        RECT 79.320 128.750 79.580 129.010 ;
        RECT 100.235 128.750 100.495 129.010 ;
        RECT 100.555 128.750 100.815 129.010 ;
        RECT 100.875 128.750 101.135 129.010 ;
        RECT 101.195 128.750 101.455 129.010 ;
        RECT 101.515 128.750 101.775 129.010 ;
        RECT 122.430 128.750 122.690 129.010 ;
        RECT 122.750 128.750 123.010 129.010 ;
        RECT 123.070 128.750 123.330 129.010 ;
        RECT 123.390 128.750 123.650 129.010 ;
        RECT 123.710 128.750 123.970 129.010 ;
        RECT 55.845 123.310 56.105 123.570 ;
        RECT 56.165 123.310 56.425 123.570 ;
        RECT 56.485 123.310 56.745 123.570 ;
        RECT 56.805 123.310 57.065 123.570 ;
        RECT 57.125 123.310 57.385 123.570 ;
        RECT 78.040 123.310 78.300 123.570 ;
        RECT 78.360 123.310 78.620 123.570 ;
        RECT 78.680 123.310 78.940 123.570 ;
        RECT 79.000 123.310 79.260 123.570 ;
        RECT 79.320 123.310 79.580 123.570 ;
        RECT 100.235 123.310 100.495 123.570 ;
        RECT 100.555 123.310 100.815 123.570 ;
        RECT 100.875 123.310 101.135 123.570 ;
        RECT 101.195 123.310 101.455 123.570 ;
        RECT 101.515 123.310 101.775 123.570 ;
        RECT 122.430 123.310 122.690 123.570 ;
        RECT 122.750 123.310 123.010 123.570 ;
        RECT 123.070 123.310 123.330 123.570 ;
        RECT 123.390 123.310 123.650 123.570 ;
        RECT 123.710 123.310 123.970 123.570 ;
        RECT 55.845 117.870 56.105 118.130 ;
        RECT 56.165 117.870 56.425 118.130 ;
        RECT 56.485 117.870 56.745 118.130 ;
        RECT 56.805 117.870 57.065 118.130 ;
        RECT 57.125 117.870 57.385 118.130 ;
        RECT 78.040 117.870 78.300 118.130 ;
        RECT 78.360 117.870 78.620 118.130 ;
        RECT 78.680 117.870 78.940 118.130 ;
        RECT 79.000 117.870 79.260 118.130 ;
        RECT 79.320 117.870 79.580 118.130 ;
        RECT 100.235 117.870 100.495 118.130 ;
        RECT 100.555 117.870 100.815 118.130 ;
        RECT 100.875 117.870 101.135 118.130 ;
        RECT 101.195 117.870 101.455 118.130 ;
        RECT 101.515 117.870 101.775 118.130 ;
        RECT 122.430 117.870 122.690 118.130 ;
        RECT 122.750 117.870 123.010 118.130 ;
        RECT 123.070 117.870 123.330 118.130 ;
        RECT 123.390 117.870 123.650 118.130 ;
        RECT 123.710 117.870 123.970 118.130 ;
        RECT 55.845 112.430 56.105 112.690 ;
        RECT 56.165 112.430 56.425 112.690 ;
        RECT 56.485 112.430 56.745 112.690 ;
        RECT 56.805 112.430 57.065 112.690 ;
        RECT 57.125 112.430 57.385 112.690 ;
        RECT 78.040 112.430 78.300 112.690 ;
        RECT 78.360 112.430 78.620 112.690 ;
        RECT 78.680 112.430 78.940 112.690 ;
        RECT 79.000 112.430 79.260 112.690 ;
        RECT 79.320 112.430 79.580 112.690 ;
        RECT 100.235 112.430 100.495 112.690 ;
        RECT 100.555 112.430 100.815 112.690 ;
        RECT 100.875 112.430 101.135 112.690 ;
        RECT 101.195 112.430 101.455 112.690 ;
        RECT 101.515 112.430 101.775 112.690 ;
        RECT 122.430 112.430 122.690 112.690 ;
        RECT 122.750 112.430 123.010 112.690 ;
        RECT 123.070 112.430 123.330 112.690 ;
        RECT 123.390 112.430 123.650 112.690 ;
        RECT 123.710 112.430 123.970 112.690 ;
        RECT 55.845 106.990 56.105 107.250 ;
        RECT 56.165 106.990 56.425 107.250 ;
        RECT 56.485 106.990 56.745 107.250 ;
        RECT 56.805 106.990 57.065 107.250 ;
        RECT 57.125 106.990 57.385 107.250 ;
        RECT 78.040 106.990 78.300 107.250 ;
        RECT 78.360 106.990 78.620 107.250 ;
        RECT 78.680 106.990 78.940 107.250 ;
        RECT 79.000 106.990 79.260 107.250 ;
        RECT 79.320 106.990 79.580 107.250 ;
        RECT 100.235 106.990 100.495 107.250 ;
        RECT 100.555 106.990 100.815 107.250 ;
        RECT 100.875 106.990 101.135 107.250 ;
        RECT 101.195 106.990 101.455 107.250 ;
        RECT 101.515 106.990 101.775 107.250 ;
        RECT 122.430 106.990 122.690 107.250 ;
        RECT 122.750 106.990 123.010 107.250 ;
        RECT 123.070 106.990 123.330 107.250 ;
        RECT 123.390 106.990 123.650 107.250 ;
        RECT 123.710 106.990 123.970 107.250 ;
        RECT 55.845 101.550 56.105 101.810 ;
        RECT 56.165 101.550 56.425 101.810 ;
        RECT 56.485 101.550 56.745 101.810 ;
        RECT 56.805 101.550 57.065 101.810 ;
        RECT 57.125 101.550 57.385 101.810 ;
        RECT 78.040 101.550 78.300 101.810 ;
        RECT 78.360 101.550 78.620 101.810 ;
        RECT 78.680 101.550 78.940 101.810 ;
        RECT 79.000 101.550 79.260 101.810 ;
        RECT 79.320 101.550 79.580 101.810 ;
        RECT 100.235 101.550 100.495 101.810 ;
        RECT 100.555 101.550 100.815 101.810 ;
        RECT 100.875 101.550 101.135 101.810 ;
        RECT 101.195 101.550 101.455 101.810 ;
        RECT 101.515 101.550 101.775 101.810 ;
        RECT 122.430 101.550 122.690 101.810 ;
        RECT 122.750 101.550 123.010 101.810 ;
        RECT 123.070 101.550 123.330 101.810 ;
        RECT 123.390 101.550 123.650 101.810 ;
        RECT 123.710 101.550 123.970 101.810 ;
        RECT 55.845 96.110 56.105 96.370 ;
        RECT 56.165 96.110 56.425 96.370 ;
        RECT 56.485 96.110 56.745 96.370 ;
        RECT 56.805 96.110 57.065 96.370 ;
        RECT 57.125 96.110 57.385 96.370 ;
        RECT 78.040 96.110 78.300 96.370 ;
        RECT 78.360 96.110 78.620 96.370 ;
        RECT 78.680 96.110 78.940 96.370 ;
        RECT 79.000 96.110 79.260 96.370 ;
        RECT 79.320 96.110 79.580 96.370 ;
        RECT 100.235 96.110 100.495 96.370 ;
        RECT 100.555 96.110 100.815 96.370 ;
        RECT 100.875 96.110 101.135 96.370 ;
        RECT 101.195 96.110 101.455 96.370 ;
        RECT 101.515 96.110 101.775 96.370 ;
        RECT 122.430 96.110 122.690 96.370 ;
        RECT 122.750 96.110 123.010 96.370 ;
        RECT 123.070 96.110 123.330 96.370 ;
        RECT 123.390 96.110 123.650 96.370 ;
        RECT 123.710 96.110 123.970 96.370 ;
        RECT 55.845 90.670 56.105 90.930 ;
        RECT 56.165 90.670 56.425 90.930 ;
        RECT 56.485 90.670 56.745 90.930 ;
        RECT 56.805 90.670 57.065 90.930 ;
        RECT 57.125 90.670 57.385 90.930 ;
        RECT 78.040 90.670 78.300 90.930 ;
        RECT 78.360 90.670 78.620 90.930 ;
        RECT 78.680 90.670 78.940 90.930 ;
        RECT 79.000 90.670 79.260 90.930 ;
        RECT 79.320 90.670 79.580 90.930 ;
        RECT 100.235 90.670 100.495 90.930 ;
        RECT 100.555 90.670 100.815 90.930 ;
        RECT 100.875 90.670 101.135 90.930 ;
        RECT 101.195 90.670 101.455 90.930 ;
        RECT 101.515 90.670 101.775 90.930 ;
        RECT 122.430 90.670 122.690 90.930 ;
        RECT 122.750 90.670 123.010 90.930 ;
        RECT 123.070 90.670 123.330 90.930 ;
        RECT 123.390 90.670 123.650 90.930 ;
        RECT 123.710 90.670 123.970 90.930 ;
        RECT 55.845 85.230 56.105 85.490 ;
        RECT 56.165 85.230 56.425 85.490 ;
        RECT 56.485 85.230 56.745 85.490 ;
        RECT 56.805 85.230 57.065 85.490 ;
        RECT 57.125 85.230 57.385 85.490 ;
        RECT 78.040 85.230 78.300 85.490 ;
        RECT 78.360 85.230 78.620 85.490 ;
        RECT 78.680 85.230 78.940 85.490 ;
        RECT 79.000 85.230 79.260 85.490 ;
        RECT 79.320 85.230 79.580 85.490 ;
        RECT 100.235 85.230 100.495 85.490 ;
        RECT 100.555 85.230 100.815 85.490 ;
        RECT 100.875 85.230 101.135 85.490 ;
        RECT 101.195 85.230 101.455 85.490 ;
        RECT 101.515 85.230 101.775 85.490 ;
        RECT 122.430 85.230 122.690 85.490 ;
        RECT 122.750 85.230 123.010 85.490 ;
        RECT 123.070 85.230 123.330 85.490 ;
        RECT 123.390 85.230 123.650 85.490 ;
        RECT 123.710 85.230 123.970 85.490 ;
        RECT 55.845 79.790 56.105 80.050 ;
        RECT 56.165 79.790 56.425 80.050 ;
        RECT 56.485 79.790 56.745 80.050 ;
        RECT 56.805 79.790 57.065 80.050 ;
        RECT 57.125 79.790 57.385 80.050 ;
        RECT 78.040 79.790 78.300 80.050 ;
        RECT 78.360 79.790 78.620 80.050 ;
        RECT 78.680 79.790 78.940 80.050 ;
        RECT 79.000 79.790 79.260 80.050 ;
        RECT 79.320 79.790 79.580 80.050 ;
        RECT 100.235 79.790 100.495 80.050 ;
        RECT 100.555 79.790 100.815 80.050 ;
        RECT 100.875 79.790 101.135 80.050 ;
        RECT 101.195 79.790 101.455 80.050 ;
        RECT 101.515 79.790 101.775 80.050 ;
        RECT 122.430 79.790 122.690 80.050 ;
        RECT 122.750 79.790 123.010 80.050 ;
        RECT 123.070 79.790 123.330 80.050 ;
        RECT 123.390 79.790 123.650 80.050 ;
        RECT 123.710 79.790 123.970 80.050 ;
        RECT 55.845 74.350 56.105 74.610 ;
        RECT 56.165 74.350 56.425 74.610 ;
        RECT 56.485 74.350 56.745 74.610 ;
        RECT 56.805 74.350 57.065 74.610 ;
        RECT 57.125 74.350 57.385 74.610 ;
        RECT 78.040 74.350 78.300 74.610 ;
        RECT 78.360 74.350 78.620 74.610 ;
        RECT 78.680 74.350 78.940 74.610 ;
        RECT 79.000 74.350 79.260 74.610 ;
        RECT 79.320 74.350 79.580 74.610 ;
        RECT 100.235 74.350 100.495 74.610 ;
        RECT 100.555 74.350 100.815 74.610 ;
        RECT 100.875 74.350 101.135 74.610 ;
        RECT 101.195 74.350 101.455 74.610 ;
        RECT 101.515 74.350 101.775 74.610 ;
        RECT 122.430 74.350 122.690 74.610 ;
        RECT 122.750 74.350 123.010 74.610 ;
        RECT 123.070 74.350 123.330 74.610 ;
        RECT 123.390 74.350 123.650 74.610 ;
        RECT 123.710 74.350 123.970 74.610 ;
        RECT 55.845 68.910 56.105 69.170 ;
        RECT 56.165 68.910 56.425 69.170 ;
        RECT 56.485 68.910 56.745 69.170 ;
        RECT 56.805 68.910 57.065 69.170 ;
        RECT 57.125 68.910 57.385 69.170 ;
        RECT 78.040 68.910 78.300 69.170 ;
        RECT 78.360 68.910 78.620 69.170 ;
        RECT 78.680 68.910 78.940 69.170 ;
        RECT 79.000 68.910 79.260 69.170 ;
        RECT 79.320 68.910 79.580 69.170 ;
        RECT 100.235 68.910 100.495 69.170 ;
        RECT 100.555 68.910 100.815 69.170 ;
        RECT 100.875 68.910 101.135 69.170 ;
        RECT 101.195 68.910 101.455 69.170 ;
        RECT 101.515 68.910 101.775 69.170 ;
        RECT 122.430 68.910 122.690 69.170 ;
        RECT 122.750 68.910 123.010 69.170 ;
        RECT 123.070 68.910 123.330 69.170 ;
        RECT 123.390 68.910 123.650 69.170 ;
        RECT 123.710 68.910 123.970 69.170 ;
        RECT 55.845 63.470 56.105 63.730 ;
        RECT 56.165 63.470 56.425 63.730 ;
        RECT 56.485 63.470 56.745 63.730 ;
        RECT 56.805 63.470 57.065 63.730 ;
        RECT 57.125 63.470 57.385 63.730 ;
        RECT 78.040 63.470 78.300 63.730 ;
        RECT 78.360 63.470 78.620 63.730 ;
        RECT 78.680 63.470 78.940 63.730 ;
        RECT 79.000 63.470 79.260 63.730 ;
        RECT 79.320 63.470 79.580 63.730 ;
        RECT 100.235 63.470 100.495 63.730 ;
        RECT 100.555 63.470 100.815 63.730 ;
        RECT 100.875 63.470 101.135 63.730 ;
        RECT 101.195 63.470 101.455 63.730 ;
        RECT 101.515 63.470 101.775 63.730 ;
        RECT 122.430 63.470 122.690 63.730 ;
        RECT 122.750 63.470 123.010 63.730 ;
        RECT 123.070 63.470 123.330 63.730 ;
        RECT 123.390 63.470 123.650 63.730 ;
        RECT 123.710 63.470 123.970 63.730 ;
      LAYER met2 ;
        RECT 55.845 134.135 57.385 134.505 ;
        RECT 78.040 134.135 79.580 134.505 ;
        RECT 100.235 134.135 101.775 134.505 ;
        RECT 122.430 134.135 123.970 134.505 ;
        RECT 55.845 128.695 57.385 129.065 ;
        RECT 78.040 128.695 79.580 129.065 ;
        RECT 100.235 128.695 101.775 129.065 ;
        RECT 122.430 128.695 123.970 129.065 ;
        RECT 55.845 123.255 57.385 123.625 ;
        RECT 78.040 123.255 79.580 123.625 ;
        RECT 100.235 123.255 101.775 123.625 ;
        RECT 122.430 123.255 123.970 123.625 ;
        RECT 55.845 117.815 57.385 118.185 ;
        RECT 78.040 117.815 79.580 118.185 ;
        RECT 100.235 117.815 101.775 118.185 ;
        RECT 122.430 117.815 123.970 118.185 ;
        RECT 55.845 112.375 57.385 112.745 ;
        RECT 78.040 112.375 79.580 112.745 ;
        RECT 100.235 112.375 101.775 112.745 ;
        RECT 122.430 112.375 123.970 112.745 ;
        RECT 55.845 106.935 57.385 107.305 ;
        RECT 78.040 106.935 79.580 107.305 ;
        RECT 100.235 106.935 101.775 107.305 ;
        RECT 122.430 106.935 123.970 107.305 ;
        RECT 55.845 101.495 57.385 101.865 ;
        RECT 78.040 101.495 79.580 101.865 ;
        RECT 100.235 101.495 101.775 101.865 ;
        RECT 122.430 101.495 123.970 101.865 ;
        RECT 55.845 96.055 57.385 96.425 ;
        RECT 78.040 96.055 79.580 96.425 ;
        RECT 100.235 96.055 101.775 96.425 ;
        RECT 122.430 96.055 123.970 96.425 ;
        RECT 55.845 90.615 57.385 90.985 ;
        RECT 78.040 90.615 79.580 90.985 ;
        RECT 100.235 90.615 101.775 90.985 ;
        RECT 122.430 90.615 123.970 90.985 ;
        RECT 55.845 85.175 57.385 85.545 ;
        RECT 78.040 85.175 79.580 85.545 ;
        RECT 100.235 85.175 101.775 85.545 ;
        RECT 122.430 85.175 123.970 85.545 ;
        RECT 55.845 79.735 57.385 80.105 ;
        RECT 78.040 79.735 79.580 80.105 ;
        RECT 100.235 79.735 101.775 80.105 ;
        RECT 122.430 79.735 123.970 80.105 ;
        RECT 55.845 74.295 57.385 74.665 ;
        RECT 78.040 74.295 79.580 74.665 ;
        RECT 100.235 74.295 101.775 74.665 ;
        RECT 122.430 74.295 123.970 74.665 ;
        RECT 55.845 68.855 57.385 69.225 ;
        RECT 78.040 68.855 79.580 69.225 ;
        RECT 100.235 68.855 101.775 69.225 ;
        RECT 122.430 68.855 123.970 69.225 ;
        RECT 55.845 63.415 57.385 63.785 ;
        RECT 78.040 63.415 79.580 63.785 ;
        RECT 100.235 63.415 101.775 63.785 ;
        RECT 122.430 63.415 123.970 63.785 ;
      LAYER via2 ;
        RECT 55.875 134.180 56.155 134.460 ;
        RECT 56.275 134.180 56.555 134.460 ;
        RECT 56.675 134.180 56.955 134.460 ;
        RECT 57.075 134.180 57.355 134.460 ;
        RECT 78.070 134.180 78.350 134.460 ;
        RECT 78.470 134.180 78.750 134.460 ;
        RECT 78.870 134.180 79.150 134.460 ;
        RECT 79.270 134.180 79.550 134.460 ;
        RECT 100.265 134.180 100.545 134.460 ;
        RECT 100.665 134.180 100.945 134.460 ;
        RECT 101.065 134.180 101.345 134.460 ;
        RECT 101.465 134.180 101.745 134.460 ;
        RECT 122.460 134.180 122.740 134.460 ;
        RECT 122.860 134.180 123.140 134.460 ;
        RECT 123.260 134.180 123.540 134.460 ;
        RECT 123.660 134.180 123.940 134.460 ;
        RECT 55.875 128.740 56.155 129.020 ;
        RECT 56.275 128.740 56.555 129.020 ;
        RECT 56.675 128.740 56.955 129.020 ;
        RECT 57.075 128.740 57.355 129.020 ;
        RECT 78.070 128.740 78.350 129.020 ;
        RECT 78.470 128.740 78.750 129.020 ;
        RECT 78.870 128.740 79.150 129.020 ;
        RECT 79.270 128.740 79.550 129.020 ;
        RECT 100.265 128.740 100.545 129.020 ;
        RECT 100.665 128.740 100.945 129.020 ;
        RECT 101.065 128.740 101.345 129.020 ;
        RECT 101.465 128.740 101.745 129.020 ;
        RECT 122.460 128.740 122.740 129.020 ;
        RECT 122.860 128.740 123.140 129.020 ;
        RECT 123.260 128.740 123.540 129.020 ;
        RECT 123.660 128.740 123.940 129.020 ;
        RECT 55.875 123.300 56.155 123.580 ;
        RECT 56.275 123.300 56.555 123.580 ;
        RECT 56.675 123.300 56.955 123.580 ;
        RECT 57.075 123.300 57.355 123.580 ;
        RECT 78.070 123.300 78.350 123.580 ;
        RECT 78.470 123.300 78.750 123.580 ;
        RECT 78.870 123.300 79.150 123.580 ;
        RECT 79.270 123.300 79.550 123.580 ;
        RECT 100.265 123.300 100.545 123.580 ;
        RECT 100.665 123.300 100.945 123.580 ;
        RECT 101.065 123.300 101.345 123.580 ;
        RECT 101.465 123.300 101.745 123.580 ;
        RECT 122.460 123.300 122.740 123.580 ;
        RECT 122.860 123.300 123.140 123.580 ;
        RECT 123.260 123.300 123.540 123.580 ;
        RECT 123.660 123.300 123.940 123.580 ;
        RECT 55.875 117.860 56.155 118.140 ;
        RECT 56.275 117.860 56.555 118.140 ;
        RECT 56.675 117.860 56.955 118.140 ;
        RECT 57.075 117.860 57.355 118.140 ;
        RECT 78.070 117.860 78.350 118.140 ;
        RECT 78.470 117.860 78.750 118.140 ;
        RECT 78.870 117.860 79.150 118.140 ;
        RECT 79.270 117.860 79.550 118.140 ;
        RECT 100.265 117.860 100.545 118.140 ;
        RECT 100.665 117.860 100.945 118.140 ;
        RECT 101.065 117.860 101.345 118.140 ;
        RECT 101.465 117.860 101.745 118.140 ;
        RECT 122.460 117.860 122.740 118.140 ;
        RECT 122.860 117.860 123.140 118.140 ;
        RECT 123.260 117.860 123.540 118.140 ;
        RECT 123.660 117.860 123.940 118.140 ;
        RECT 55.875 112.420 56.155 112.700 ;
        RECT 56.275 112.420 56.555 112.700 ;
        RECT 56.675 112.420 56.955 112.700 ;
        RECT 57.075 112.420 57.355 112.700 ;
        RECT 78.070 112.420 78.350 112.700 ;
        RECT 78.470 112.420 78.750 112.700 ;
        RECT 78.870 112.420 79.150 112.700 ;
        RECT 79.270 112.420 79.550 112.700 ;
        RECT 100.265 112.420 100.545 112.700 ;
        RECT 100.665 112.420 100.945 112.700 ;
        RECT 101.065 112.420 101.345 112.700 ;
        RECT 101.465 112.420 101.745 112.700 ;
        RECT 122.460 112.420 122.740 112.700 ;
        RECT 122.860 112.420 123.140 112.700 ;
        RECT 123.260 112.420 123.540 112.700 ;
        RECT 123.660 112.420 123.940 112.700 ;
        RECT 55.875 106.980 56.155 107.260 ;
        RECT 56.275 106.980 56.555 107.260 ;
        RECT 56.675 106.980 56.955 107.260 ;
        RECT 57.075 106.980 57.355 107.260 ;
        RECT 78.070 106.980 78.350 107.260 ;
        RECT 78.470 106.980 78.750 107.260 ;
        RECT 78.870 106.980 79.150 107.260 ;
        RECT 79.270 106.980 79.550 107.260 ;
        RECT 100.265 106.980 100.545 107.260 ;
        RECT 100.665 106.980 100.945 107.260 ;
        RECT 101.065 106.980 101.345 107.260 ;
        RECT 101.465 106.980 101.745 107.260 ;
        RECT 122.460 106.980 122.740 107.260 ;
        RECT 122.860 106.980 123.140 107.260 ;
        RECT 123.260 106.980 123.540 107.260 ;
        RECT 123.660 106.980 123.940 107.260 ;
        RECT 55.875 101.540 56.155 101.820 ;
        RECT 56.275 101.540 56.555 101.820 ;
        RECT 56.675 101.540 56.955 101.820 ;
        RECT 57.075 101.540 57.355 101.820 ;
        RECT 78.070 101.540 78.350 101.820 ;
        RECT 78.470 101.540 78.750 101.820 ;
        RECT 78.870 101.540 79.150 101.820 ;
        RECT 79.270 101.540 79.550 101.820 ;
        RECT 100.265 101.540 100.545 101.820 ;
        RECT 100.665 101.540 100.945 101.820 ;
        RECT 101.065 101.540 101.345 101.820 ;
        RECT 101.465 101.540 101.745 101.820 ;
        RECT 122.460 101.540 122.740 101.820 ;
        RECT 122.860 101.540 123.140 101.820 ;
        RECT 123.260 101.540 123.540 101.820 ;
        RECT 123.660 101.540 123.940 101.820 ;
        RECT 55.875 96.100 56.155 96.380 ;
        RECT 56.275 96.100 56.555 96.380 ;
        RECT 56.675 96.100 56.955 96.380 ;
        RECT 57.075 96.100 57.355 96.380 ;
        RECT 78.070 96.100 78.350 96.380 ;
        RECT 78.470 96.100 78.750 96.380 ;
        RECT 78.870 96.100 79.150 96.380 ;
        RECT 79.270 96.100 79.550 96.380 ;
        RECT 100.265 96.100 100.545 96.380 ;
        RECT 100.665 96.100 100.945 96.380 ;
        RECT 101.065 96.100 101.345 96.380 ;
        RECT 101.465 96.100 101.745 96.380 ;
        RECT 122.460 96.100 122.740 96.380 ;
        RECT 122.860 96.100 123.140 96.380 ;
        RECT 123.260 96.100 123.540 96.380 ;
        RECT 123.660 96.100 123.940 96.380 ;
        RECT 55.875 90.660 56.155 90.940 ;
        RECT 56.275 90.660 56.555 90.940 ;
        RECT 56.675 90.660 56.955 90.940 ;
        RECT 57.075 90.660 57.355 90.940 ;
        RECT 78.070 90.660 78.350 90.940 ;
        RECT 78.470 90.660 78.750 90.940 ;
        RECT 78.870 90.660 79.150 90.940 ;
        RECT 79.270 90.660 79.550 90.940 ;
        RECT 100.265 90.660 100.545 90.940 ;
        RECT 100.665 90.660 100.945 90.940 ;
        RECT 101.065 90.660 101.345 90.940 ;
        RECT 101.465 90.660 101.745 90.940 ;
        RECT 122.460 90.660 122.740 90.940 ;
        RECT 122.860 90.660 123.140 90.940 ;
        RECT 123.260 90.660 123.540 90.940 ;
        RECT 123.660 90.660 123.940 90.940 ;
        RECT 55.875 85.220 56.155 85.500 ;
        RECT 56.275 85.220 56.555 85.500 ;
        RECT 56.675 85.220 56.955 85.500 ;
        RECT 57.075 85.220 57.355 85.500 ;
        RECT 78.070 85.220 78.350 85.500 ;
        RECT 78.470 85.220 78.750 85.500 ;
        RECT 78.870 85.220 79.150 85.500 ;
        RECT 79.270 85.220 79.550 85.500 ;
        RECT 100.265 85.220 100.545 85.500 ;
        RECT 100.665 85.220 100.945 85.500 ;
        RECT 101.065 85.220 101.345 85.500 ;
        RECT 101.465 85.220 101.745 85.500 ;
        RECT 122.460 85.220 122.740 85.500 ;
        RECT 122.860 85.220 123.140 85.500 ;
        RECT 123.260 85.220 123.540 85.500 ;
        RECT 123.660 85.220 123.940 85.500 ;
        RECT 55.875 79.780 56.155 80.060 ;
        RECT 56.275 79.780 56.555 80.060 ;
        RECT 56.675 79.780 56.955 80.060 ;
        RECT 57.075 79.780 57.355 80.060 ;
        RECT 78.070 79.780 78.350 80.060 ;
        RECT 78.470 79.780 78.750 80.060 ;
        RECT 78.870 79.780 79.150 80.060 ;
        RECT 79.270 79.780 79.550 80.060 ;
        RECT 100.265 79.780 100.545 80.060 ;
        RECT 100.665 79.780 100.945 80.060 ;
        RECT 101.065 79.780 101.345 80.060 ;
        RECT 101.465 79.780 101.745 80.060 ;
        RECT 122.460 79.780 122.740 80.060 ;
        RECT 122.860 79.780 123.140 80.060 ;
        RECT 123.260 79.780 123.540 80.060 ;
        RECT 123.660 79.780 123.940 80.060 ;
        RECT 55.875 74.340 56.155 74.620 ;
        RECT 56.275 74.340 56.555 74.620 ;
        RECT 56.675 74.340 56.955 74.620 ;
        RECT 57.075 74.340 57.355 74.620 ;
        RECT 78.070 74.340 78.350 74.620 ;
        RECT 78.470 74.340 78.750 74.620 ;
        RECT 78.870 74.340 79.150 74.620 ;
        RECT 79.270 74.340 79.550 74.620 ;
        RECT 100.265 74.340 100.545 74.620 ;
        RECT 100.665 74.340 100.945 74.620 ;
        RECT 101.065 74.340 101.345 74.620 ;
        RECT 101.465 74.340 101.745 74.620 ;
        RECT 122.460 74.340 122.740 74.620 ;
        RECT 122.860 74.340 123.140 74.620 ;
        RECT 123.260 74.340 123.540 74.620 ;
        RECT 123.660 74.340 123.940 74.620 ;
        RECT 55.875 68.900 56.155 69.180 ;
        RECT 56.275 68.900 56.555 69.180 ;
        RECT 56.675 68.900 56.955 69.180 ;
        RECT 57.075 68.900 57.355 69.180 ;
        RECT 78.070 68.900 78.350 69.180 ;
        RECT 78.470 68.900 78.750 69.180 ;
        RECT 78.870 68.900 79.150 69.180 ;
        RECT 79.270 68.900 79.550 69.180 ;
        RECT 100.265 68.900 100.545 69.180 ;
        RECT 100.665 68.900 100.945 69.180 ;
        RECT 101.065 68.900 101.345 69.180 ;
        RECT 101.465 68.900 101.745 69.180 ;
        RECT 122.460 68.900 122.740 69.180 ;
        RECT 122.860 68.900 123.140 69.180 ;
        RECT 123.260 68.900 123.540 69.180 ;
        RECT 123.660 68.900 123.940 69.180 ;
        RECT 55.875 63.460 56.155 63.740 ;
        RECT 56.275 63.460 56.555 63.740 ;
        RECT 56.675 63.460 56.955 63.740 ;
        RECT 57.075 63.460 57.355 63.740 ;
        RECT 78.070 63.460 78.350 63.740 ;
        RECT 78.470 63.460 78.750 63.740 ;
        RECT 78.870 63.460 79.150 63.740 ;
        RECT 79.270 63.460 79.550 63.740 ;
        RECT 100.265 63.460 100.545 63.740 ;
        RECT 100.665 63.460 100.945 63.740 ;
        RECT 101.065 63.460 101.345 63.740 ;
        RECT 101.465 63.460 101.745 63.740 ;
        RECT 122.460 63.460 122.740 63.740 ;
        RECT 122.860 63.460 123.140 63.740 ;
        RECT 123.260 63.460 123.540 63.740 ;
        RECT 123.660 63.460 123.940 63.740 ;
      LAYER met3 ;
        RECT 55.825 134.155 57.405 134.485 ;
        RECT 78.020 134.155 79.600 134.485 ;
        RECT 100.215 134.155 101.795 134.485 ;
        RECT 122.410 134.155 123.990 134.485 ;
        RECT 55.825 128.715 57.405 129.045 ;
        RECT 78.020 128.715 79.600 129.045 ;
        RECT 100.215 128.715 101.795 129.045 ;
        RECT 122.410 128.715 123.990 129.045 ;
        RECT 55.825 123.275 57.405 123.605 ;
        RECT 78.020 123.275 79.600 123.605 ;
        RECT 100.215 123.275 101.795 123.605 ;
        RECT 122.410 123.275 123.990 123.605 ;
        RECT 55.825 117.835 57.405 118.165 ;
        RECT 78.020 117.835 79.600 118.165 ;
        RECT 100.215 117.835 101.795 118.165 ;
        RECT 122.410 117.835 123.990 118.165 ;
        RECT 55.825 112.395 57.405 112.725 ;
        RECT 78.020 112.395 79.600 112.725 ;
        RECT 100.215 112.395 101.795 112.725 ;
        RECT 122.410 112.395 123.990 112.725 ;
        RECT 55.825 106.955 57.405 107.285 ;
        RECT 78.020 106.955 79.600 107.285 ;
        RECT 100.215 106.955 101.795 107.285 ;
        RECT 122.410 106.955 123.990 107.285 ;
        RECT 55.825 101.515 57.405 101.845 ;
        RECT 78.020 101.515 79.600 101.845 ;
        RECT 100.215 101.515 101.795 101.845 ;
        RECT 122.410 101.515 123.990 101.845 ;
        RECT 55.825 96.075 57.405 96.405 ;
        RECT 78.020 96.075 79.600 96.405 ;
        RECT 100.215 96.075 101.795 96.405 ;
        RECT 122.410 96.075 123.990 96.405 ;
        RECT 55.825 90.635 57.405 90.965 ;
        RECT 78.020 90.635 79.600 90.965 ;
        RECT 100.215 90.635 101.795 90.965 ;
        RECT 122.410 90.635 123.990 90.965 ;
        RECT 55.825 85.195 57.405 85.525 ;
        RECT 78.020 85.195 79.600 85.525 ;
        RECT 100.215 85.195 101.795 85.525 ;
        RECT 122.410 85.195 123.990 85.525 ;
        RECT 55.825 79.755 57.405 80.085 ;
        RECT 78.020 79.755 79.600 80.085 ;
        RECT 100.215 79.755 101.795 80.085 ;
        RECT 122.410 79.755 123.990 80.085 ;
        RECT 55.825 74.315 57.405 74.645 ;
        RECT 78.020 74.315 79.600 74.645 ;
        RECT 100.215 74.315 101.795 74.645 ;
        RECT 122.410 74.315 123.990 74.645 ;
        RECT 55.825 68.875 57.405 69.205 ;
        RECT 78.020 68.875 79.600 69.205 ;
        RECT 100.215 68.875 101.795 69.205 ;
        RECT 122.410 68.875 123.990 69.205 ;
        RECT 55.825 63.435 57.405 63.765 ;
        RECT 78.020 63.435 79.600 63.765 ;
        RECT 100.215 63.435 101.795 63.765 ;
        RECT 122.410 63.435 123.990 63.765 ;
      LAYER via3 ;
        RECT 55.855 134.160 56.175 134.480 ;
        RECT 56.255 134.160 56.575 134.480 ;
        RECT 56.655 134.160 56.975 134.480 ;
        RECT 57.055 134.160 57.375 134.480 ;
        RECT 78.050 134.160 78.370 134.480 ;
        RECT 78.450 134.160 78.770 134.480 ;
        RECT 78.850 134.160 79.170 134.480 ;
        RECT 79.250 134.160 79.570 134.480 ;
        RECT 100.245 134.160 100.565 134.480 ;
        RECT 100.645 134.160 100.965 134.480 ;
        RECT 101.045 134.160 101.365 134.480 ;
        RECT 101.445 134.160 101.765 134.480 ;
        RECT 122.440 134.160 122.760 134.480 ;
        RECT 122.840 134.160 123.160 134.480 ;
        RECT 123.240 134.160 123.560 134.480 ;
        RECT 123.640 134.160 123.960 134.480 ;
        RECT 55.855 128.720 56.175 129.040 ;
        RECT 56.255 128.720 56.575 129.040 ;
        RECT 56.655 128.720 56.975 129.040 ;
        RECT 57.055 128.720 57.375 129.040 ;
        RECT 78.050 128.720 78.370 129.040 ;
        RECT 78.450 128.720 78.770 129.040 ;
        RECT 78.850 128.720 79.170 129.040 ;
        RECT 79.250 128.720 79.570 129.040 ;
        RECT 100.245 128.720 100.565 129.040 ;
        RECT 100.645 128.720 100.965 129.040 ;
        RECT 101.045 128.720 101.365 129.040 ;
        RECT 101.445 128.720 101.765 129.040 ;
        RECT 122.440 128.720 122.760 129.040 ;
        RECT 122.840 128.720 123.160 129.040 ;
        RECT 123.240 128.720 123.560 129.040 ;
        RECT 123.640 128.720 123.960 129.040 ;
        RECT 55.855 123.280 56.175 123.600 ;
        RECT 56.255 123.280 56.575 123.600 ;
        RECT 56.655 123.280 56.975 123.600 ;
        RECT 57.055 123.280 57.375 123.600 ;
        RECT 78.050 123.280 78.370 123.600 ;
        RECT 78.450 123.280 78.770 123.600 ;
        RECT 78.850 123.280 79.170 123.600 ;
        RECT 79.250 123.280 79.570 123.600 ;
        RECT 100.245 123.280 100.565 123.600 ;
        RECT 100.645 123.280 100.965 123.600 ;
        RECT 101.045 123.280 101.365 123.600 ;
        RECT 101.445 123.280 101.765 123.600 ;
        RECT 122.440 123.280 122.760 123.600 ;
        RECT 122.840 123.280 123.160 123.600 ;
        RECT 123.240 123.280 123.560 123.600 ;
        RECT 123.640 123.280 123.960 123.600 ;
        RECT 55.855 117.840 56.175 118.160 ;
        RECT 56.255 117.840 56.575 118.160 ;
        RECT 56.655 117.840 56.975 118.160 ;
        RECT 57.055 117.840 57.375 118.160 ;
        RECT 78.050 117.840 78.370 118.160 ;
        RECT 78.450 117.840 78.770 118.160 ;
        RECT 78.850 117.840 79.170 118.160 ;
        RECT 79.250 117.840 79.570 118.160 ;
        RECT 100.245 117.840 100.565 118.160 ;
        RECT 100.645 117.840 100.965 118.160 ;
        RECT 101.045 117.840 101.365 118.160 ;
        RECT 101.445 117.840 101.765 118.160 ;
        RECT 122.440 117.840 122.760 118.160 ;
        RECT 122.840 117.840 123.160 118.160 ;
        RECT 123.240 117.840 123.560 118.160 ;
        RECT 123.640 117.840 123.960 118.160 ;
        RECT 55.855 112.400 56.175 112.720 ;
        RECT 56.255 112.400 56.575 112.720 ;
        RECT 56.655 112.400 56.975 112.720 ;
        RECT 57.055 112.400 57.375 112.720 ;
        RECT 78.050 112.400 78.370 112.720 ;
        RECT 78.450 112.400 78.770 112.720 ;
        RECT 78.850 112.400 79.170 112.720 ;
        RECT 79.250 112.400 79.570 112.720 ;
        RECT 100.245 112.400 100.565 112.720 ;
        RECT 100.645 112.400 100.965 112.720 ;
        RECT 101.045 112.400 101.365 112.720 ;
        RECT 101.445 112.400 101.765 112.720 ;
        RECT 122.440 112.400 122.760 112.720 ;
        RECT 122.840 112.400 123.160 112.720 ;
        RECT 123.240 112.400 123.560 112.720 ;
        RECT 123.640 112.400 123.960 112.720 ;
        RECT 55.855 106.960 56.175 107.280 ;
        RECT 56.255 106.960 56.575 107.280 ;
        RECT 56.655 106.960 56.975 107.280 ;
        RECT 57.055 106.960 57.375 107.280 ;
        RECT 78.050 106.960 78.370 107.280 ;
        RECT 78.450 106.960 78.770 107.280 ;
        RECT 78.850 106.960 79.170 107.280 ;
        RECT 79.250 106.960 79.570 107.280 ;
        RECT 100.245 106.960 100.565 107.280 ;
        RECT 100.645 106.960 100.965 107.280 ;
        RECT 101.045 106.960 101.365 107.280 ;
        RECT 101.445 106.960 101.765 107.280 ;
        RECT 122.440 106.960 122.760 107.280 ;
        RECT 122.840 106.960 123.160 107.280 ;
        RECT 123.240 106.960 123.560 107.280 ;
        RECT 123.640 106.960 123.960 107.280 ;
        RECT 55.855 101.520 56.175 101.840 ;
        RECT 56.255 101.520 56.575 101.840 ;
        RECT 56.655 101.520 56.975 101.840 ;
        RECT 57.055 101.520 57.375 101.840 ;
        RECT 78.050 101.520 78.370 101.840 ;
        RECT 78.450 101.520 78.770 101.840 ;
        RECT 78.850 101.520 79.170 101.840 ;
        RECT 79.250 101.520 79.570 101.840 ;
        RECT 100.245 101.520 100.565 101.840 ;
        RECT 100.645 101.520 100.965 101.840 ;
        RECT 101.045 101.520 101.365 101.840 ;
        RECT 101.445 101.520 101.765 101.840 ;
        RECT 122.440 101.520 122.760 101.840 ;
        RECT 122.840 101.520 123.160 101.840 ;
        RECT 123.240 101.520 123.560 101.840 ;
        RECT 123.640 101.520 123.960 101.840 ;
        RECT 55.855 96.080 56.175 96.400 ;
        RECT 56.255 96.080 56.575 96.400 ;
        RECT 56.655 96.080 56.975 96.400 ;
        RECT 57.055 96.080 57.375 96.400 ;
        RECT 78.050 96.080 78.370 96.400 ;
        RECT 78.450 96.080 78.770 96.400 ;
        RECT 78.850 96.080 79.170 96.400 ;
        RECT 79.250 96.080 79.570 96.400 ;
        RECT 100.245 96.080 100.565 96.400 ;
        RECT 100.645 96.080 100.965 96.400 ;
        RECT 101.045 96.080 101.365 96.400 ;
        RECT 101.445 96.080 101.765 96.400 ;
        RECT 122.440 96.080 122.760 96.400 ;
        RECT 122.840 96.080 123.160 96.400 ;
        RECT 123.240 96.080 123.560 96.400 ;
        RECT 123.640 96.080 123.960 96.400 ;
        RECT 55.855 90.640 56.175 90.960 ;
        RECT 56.255 90.640 56.575 90.960 ;
        RECT 56.655 90.640 56.975 90.960 ;
        RECT 57.055 90.640 57.375 90.960 ;
        RECT 78.050 90.640 78.370 90.960 ;
        RECT 78.450 90.640 78.770 90.960 ;
        RECT 78.850 90.640 79.170 90.960 ;
        RECT 79.250 90.640 79.570 90.960 ;
        RECT 100.245 90.640 100.565 90.960 ;
        RECT 100.645 90.640 100.965 90.960 ;
        RECT 101.045 90.640 101.365 90.960 ;
        RECT 101.445 90.640 101.765 90.960 ;
        RECT 122.440 90.640 122.760 90.960 ;
        RECT 122.840 90.640 123.160 90.960 ;
        RECT 123.240 90.640 123.560 90.960 ;
        RECT 123.640 90.640 123.960 90.960 ;
        RECT 55.855 85.200 56.175 85.520 ;
        RECT 56.255 85.200 56.575 85.520 ;
        RECT 56.655 85.200 56.975 85.520 ;
        RECT 57.055 85.200 57.375 85.520 ;
        RECT 78.050 85.200 78.370 85.520 ;
        RECT 78.450 85.200 78.770 85.520 ;
        RECT 78.850 85.200 79.170 85.520 ;
        RECT 79.250 85.200 79.570 85.520 ;
        RECT 100.245 85.200 100.565 85.520 ;
        RECT 100.645 85.200 100.965 85.520 ;
        RECT 101.045 85.200 101.365 85.520 ;
        RECT 101.445 85.200 101.765 85.520 ;
        RECT 122.440 85.200 122.760 85.520 ;
        RECT 122.840 85.200 123.160 85.520 ;
        RECT 123.240 85.200 123.560 85.520 ;
        RECT 123.640 85.200 123.960 85.520 ;
        RECT 55.855 79.760 56.175 80.080 ;
        RECT 56.255 79.760 56.575 80.080 ;
        RECT 56.655 79.760 56.975 80.080 ;
        RECT 57.055 79.760 57.375 80.080 ;
        RECT 78.050 79.760 78.370 80.080 ;
        RECT 78.450 79.760 78.770 80.080 ;
        RECT 78.850 79.760 79.170 80.080 ;
        RECT 79.250 79.760 79.570 80.080 ;
        RECT 100.245 79.760 100.565 80.080 ;
        RECT 100.645 79.760 100.965 80.080 ;
        RECT 101.045 79.760 101.365 80.080 ;
        RECT 101.445 79.760 101.765 80.080 ;
        RECT 122.440 79.760 122.760 80.080 ;
        RECT 122.840 79.760 123.160 80.080 ;
        RECT 123.240 79.760 123.560 80.080 ;
        RECT 123.640 79.760 123.960 80.080 ;
        RECT 55.855 74.320 56.175 74.640 ;
        RECT 56.255 74.320 56.575 74.640 ;
        RECT 56.655 74.320 56.975 74.640 ;
        RECT 57.055 74.320 57.375 74.640 ;
        RECT 78.050 74.320 78.370 74.640 ;
        RECT 78.450 74.320 78.770 74.640 ;
        RECT 78.850 74.320 79.170 74.640 ;
        RECT 79.250 74.320 79.570 74.640 ;
        RECT 100.245 74.320 100.565 74.640 ;
        RECT 100.645 74.320 100.965 74.640 ;
        RECT 101.045 74.320 101.365 74.640 ;
        RECT 101.445 74.320 101.765 74.640 ;
        RECT 122.440 74.320 122.760 74.640 ;
        RECT 122.840 74.320 123.160 74.640 ;
        RECT 123.240 74.320 123.560 74.640 ;
        RECT 123.640 74.320 123.960 74.640 ;
        RECT 55.855 68.880 56.175 69.200 ;
        RECT 56.255 68.880 56.575 69.200 ;
        RECT 56.655 68.880 56.975 69.200 ;
        RECT 57.055 68.880 57.375 69.200 ;
        RECT 78.050 68.880 78.370 69.200 ;
        RECT 78.450 68.880 78.770 69.200 ;
        RECT 78.850 68.880 79.170 69.200 ;
        RECT 79.250 68.880 79.570 69.200 ;
        RECT 100.245 68.880 100.565 69.200 ;
        RECT 100.645 68.880 100.965 69.200 ;
        RECT 101.045 68.880 101.365 69.200 ;
        RECT 101.445 68.880 101.765 69.200 ;
        RECT 122.440 68.880 122.760 69.200 ;
        RECT 122.840 68.880 123.160 69.200 ;
        RECT 123.240 68.880 123.560 69.200 ;
        RECT 123.640 68.880 123.960 69.200 ;
        RECT 55.855 63.440 56.175 63.760 ;
        RECT 56.255 63.440 56.575 63.760 ;
        RECT 56.655 63.440 56.975 63.760 ;
        RECT 57.055 63.440 57.375 63.760 ;
        RECT 78.050 63.440 78.370 63.760 ;
        RECT 78.450 63.440 78.770 63.760 ;
        RECT 78.850 63.440 79.170 63.760 ;
        RECT 79.250 63.440 79.570 63.760 ;
        RECT 100.245 63.440 100.565 63.760 ;
        RECT 100.645 63.440 100.965 63.760 ;
        RECT 101.045 63.440 101.365 63.760 ;
        RECT 101.445 63.440 101.765 63.760 ;
        RECT 122.440 63.440 122.760 63.760 ;
        RECT 122.840 63.440 123.160 63.760 ;
        RECT 123.240 63.440 123.560 63.760 ;
        RECT 123.640 63.440 123.960 63.760 ;
      LAYER met4 ;
        RECT 55.815 60.640 57.415 137.280 ;
        RECT 78.010 60.640 79.610 137.280 ;
        RECT 100.205 60.640 101.805 137.280 ;
        RECT 122.400 60.640 124.000 137.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 58.545 136.195 58.715 136.720 ;
        RECT 71.425 136.195 71.595 136.720 ;
        RECT 84.305 136.195 84.475 136.720 ;
        RECT 97.185 136.195 97.355 136.720 ;
        RECT 110.065 136.195 110.235 136.720 ;
        RECT 122.945 136.195 123.115 136.720 ;
        RECT 58.545 131.920 58.715 132.445 ;
        RECT 84.305 131.920 84.475 132.445 ;
        RECT 110.065 131.920 110.235 132.445 ;
        RECT 71.425 130.755 71.595 131.280 ;
        RECT 97.185 130.755 97.355 131.280 ;
        RECT 122.945 130.755 123.115 131.280 ;
        RECT 58.545 126.480 58.715 127.005 ;
        RECT 84.305 126.480 84.475 127.005 ;
        RECT 110.065 126.480 110.235 127.005 ;
        RECT 71.425 125.315 71.595 125.840 ;
        RECT 97.185 125.315 97.355 125.840 ;
        RECT 122.945 125.315 123.115 125.840 ;
        RECT 58.545 121.040 58.715 121.565 ;
        RECT 84.305 121.040 84.475 121.565 ;
        RECT 110.065 121.040 110.235 121.565 ;
        RECT 71.425 119.875 71.595 120.400 ;
        RECT 97.185 119.875 97.355 120.400 ;
        RECT 122.945 119.875 123.115 120.400 ;
        RECT 58.545 115.600 58.715 116.125 ;
        RECT 84.305 115.600 84.475 116.125 ;
        RECT 110.065 115.600 110.235 116.125 ;
        RECT 71.425 114.435 71.595 114.960 ;
        RECT 97.185 114.435 97.355 114.960 ;
        RECT 122.945 114.435 123.115 114.960 ;
        RECT 58.545 110.160 58.715 110.685 ;
        RECT 84.305 110.160 84.475 110.685 ;
        RECT 110.065 110.160 110.235 110.685 ;
        RECT 71.425 108.995 71.595 109.520 ;
        RECT 97.185 108.995 97.355 109.520 ;
        RECT 122.945 108.995 123.115 109.520 ;
        RECT 58.545 104.720 58.715 105.245 ;
        RECT 84.305 104.720 84.475 105.245 ;
        RECT 110.065 104.720 110.235 105.245 ;
        RECT 71.425 103.555 71.595 104.080 ;
        RECT 97.185 103.555 97.355 104.080 ;
        RECT 122.945 103.555 123.115 104.080 ;
        RECT 58.545 99.280 58.715 99.805 ;
        RECT 84.305 99.280 84.475 99.805 ;
        RECT 110.065 99.280 110.235 99.805 ;
        RECT 71.425 98.115 71.595 98.640 ;
        RECT 97.185 98.115 97.355 98.640 ;
        RECT 122.945 98.115 123.115 98.640 ;
        RECT 58.545 93.840 58.715 94.365 ;
        RECT 84.305 93.840 84.475 94.365 ;
        RECT 110.065 93.840 110.235 94.365 ;
        RECT 71.425 92.675 71.595 93.200 ;
        RECT 97.185 92.675 97.355 93.200 ;
        RECT 122.945 92.675 123.115 93.200 ;
        RECT 58.545 88.400 58.715 88.925 ;
        RECT 84.305 88.400 84.475 88.925 ;
        RECT 110.065 88.400 110.235 88.925 ;
        RECT 71.425 87.235 71.595 87.760 ;
        RECT 97.185 87.235 97.355 87.760 ;
        RECT 122.945 87.235 123.115 87.760 ;
        RECT 58.545 82.960 58.715 83.485 ;
        RECT 84.305 82.960 84.475 83.485 ;
        RECT 110.065 82.960 110.235 83.485 ;
        RECT 71.425 81.795 71.595 82.320 ;
        RECT 97.185 81.795 97.355 82.320 ;
        RECT 122.945 81.795 123.115 82.320 ;
        RECT 58.545 77.520 58.715 78.045 ;
        RECT 84.305 77.520 84.475 78.045 ;
        RECT 110.065 77.520 110.235 78.045 ;
        RECT 71.425 76.355 71.595 76.880 ;
        RECT 97.185 76.355 97.355 76.880 ;
        RECT 122.945 76.355 123.115 76.880 ;
        RECT 58.545 72.080 58.715 72.605 ;
        RECT 84.305 72.080 84.475 72.605 ;
        RECT 110.065 72.080 110.235 72.605 ;
        RECT 71.425 70.915 71.595 71.440 ;
        RECT 97.185 70.915 97.355 71.440 ;
        RECT 122.945 70.915 123.115 71.440 ;
        RECT 58.545 66.640 58.715 67.165 ;
        RECT 84.305 66.640 84.475 67.165 ;
        RECT 110.065 66.640 110.235 67.165 ;
        RECT 71.425 65.475 71.595 66.000 ;
        RECT 97.185 65.475 97.355 66.000 ;
        RECT 122.945 65.475 123.115 66.000 ;
        RECT 58.545 61.200 58.715 61.725 ;
        RECT 71.425 61.200 71.595 61.725 ;
        RECT 84.305 61.200 84.475 61.725 ;
        RECT 97.185 61.200 97.355 61.725 ;
        RECT 110.065 61.200 110.235 61.725 ;
        RECT 122.945 61.200 123.115 61.725 ;
      LAYER li1 ;
        RECT 45.520 136.955 134.300 137.125 ;
        RECT 45.605 136.205 46.815 136.955 ;
        RECT 46.985 136.410 52.330 136.955 ;
        RECT 52.505 136.410 57.850 136.955 ;
        RECT 45.605 135.665 46.125 136.205 ;
        RECT 48.570 135.580 48.910 136.410 ;
        RECT 54.090 135.580 54.430 136.410 ;
        RECT 58.485 136.230 58.775 136.955 ;
        RECT 58.945 136.410 64.290 136.955 ;
        RECT 64.465 136.410 69.810 136.955 ;
        RECT 60.530 135.580 60.870 136.410 ;
        RECT 66.050 135.580 66.390 136.410 ;
        RECT 69.985 136.205 71.195 136.955 ;
        RECT 71.365 136.230 71.655 136.955 ;
        RECT 71.825 136.410 77.170 136.955 ;
        RECT 77.345 136.410 82.690 136.955 ;
        RECT 69.985 135.665 70.505 136.205 ;
        RECT 73.410 135.580 73.750 136.410 ;
        RECT 78.930 135.580 79.270 136.410 ;
        RECT 82.865 136.205 84.075 136.955 ;
        RECT 84.245 136.230 84.535 136.955 ;
        RECT 84.705 136.410 90.050 136.955 ;
        RECT 90.225 136.410 95.570 136.955 ;
        RECT 82.865 135.665 83.385 136.205 ;
        RECT 86.290 135.580 86.630 136.410 ;
        RECT 91.810 135.580 92.150 136.410 ;
        RECT 95.745 136.205 96.955 136.955 ;
        RECT 97.125 136.230 97.415 136.955 ;
        RECT 97.585 136.410 102.930 136.955 ;
        RECT 103.105 136.410 108.450 136.955 ;
        RECT 95.745 135.665 96.265 136.205 ;
        RECT 99.170 135.580 99.510 136.410 ;
        RECT 104.690 135.580 105.030 136.410 ;
        RECT 108.625 136.205 109.835 136.955 ;
        RECT 110.005 136.230 110.295 136.955 ;
        RECT 110.465 136.410 115.810 136.955 ;
        RECT 115.985 136.410 121.330 136.955 ;
        RECT 108.625 135.665 109.145 136.205 ;
        RECT 112.050 135.580 112.390 136.410 ;
        RECT 117.570 135.580 117.910 136.410 ;
        RECT 121.505 136.205 122.715 136.955 ;
        RECT 122.885 136.230 123.175 136.955 ;
        RECT 123.345 136.410 128.690 136.955 ;
        RECT 121.505 135.665 122.025 136.205 ;
        RECT 124.930 135.580 125.270 136.410 ;
        RECT 128.865 136.185 132.375 136.955 ;
        RECT 133.005 136.205 134.215 136.955 ;
        RECT 128.865 135.665 130.515 136.185 ;
        RECT 133.695 135.665 134.215 136.205 ;
        RECT 45.605 132.435 46.125 132.975 ;
        RECT 45.605 131.685 46.815 132.435 ;
        RECT 48.570 132.230 48.910 133.060 ;
        RECT 54.090 132.230 54.430 133.060 ;
        RECT 46.985 131.685 52.330 132.230 ;
        RECT 52.505 131.685 57.850 132.230 ;
        RECT 58.485 131.685 58.775 132.410 ;
        RECT 60.530 132.230 60.870 133.060 ;
        RECT 66.050 132.230 66.390 133.060 ;
        RECT 71.570 132.230 71.910 133.060 ;
        RECT 77.090 132.230 77.430 133.060 ;
        RECT 81.025 132.455 82.235 132.975 ;
        RECT 58.945 131.685 64.290 132.230 ;
        RECT 64.465 131.685 69.810 132.230 ;
        RECT 69.985 131.685 75.330 132.230 ;
        RECT 75.505 131.685 80.850 132.230 ;
        RECT 81.025 131.685 83.615 132.455 ;
        RECT 84.245 131.685 84.535 132.410 ;
        RECT 86.290 132.230 86.630 133.060 ;
        RECT 91.810 132.230 92.150 133.060 ;
        RECT 97.330 132.230 97.670 133.060 ;
        RECT 102.850 132.230 103.190 133.060 ;
        RECT 106.785 132.455 107.995 132.975 ;
        RECT 84.705 131.685 90.050 132.230 ;
        RECT 90.225 131.685 95.570 132.230 ;
        RECT 95.745 131.685 101.090 132.230 ;
        RECT 101.265 131.685 106.610 132.230 ;
        RECT 106.785 131.685 109.375 132.455 ;
        RECT 110.005 131.685 110.295 132.410 ;
        RECT 112.050 132.230 112.390 133.060 ;
        RECT 117.570 132.230 117.910 133.060 ;
        RECT 123.090 132.230 123.430 133.060 ;
        RECT 128.610 132.230 128.950 133.060 ;
        RECT 133.695 132.435 134.215 132.975 ;
        RECT 110.465 131.685 115.810 132.230 ;
        RECT 115.985 131.685 121.330 132.230 ;
        RECT 121.505 131.685 126.850 132.230 ;
        RECT 127.025 131.685 132.370 132.230 ;
        RECT 133.005 131.685 134.215 132.435 ;
        RECT 45.520 131.515 134.300 131.685 ;
        RECT 45.605 130.765 46.815 131.515 ;
        RECT 46.985 130.970 52.330 131.515 ;
        RECT 52.505 130.970 57.850 131.515 ;
        RECT 58.025 130.970 63.370 131.515 ;
        RECT 63.545 130.970 68.890 131.515 ;
        RECT 45.605 130.225 46.125 130.765 ;
        RECT 48.570 130.140 48.910 130.970 ;
        RECT 54.090 130.140 54.430 130.970 ;
        RECT 59.610 130.140 59.950 130.970 ;
        RECT 65.130 130.140 65.470 130.970 ;
        RECT 69.065 130.745 70.735 131.515 ;
        RECT 71.365 130.790 71.655 131.515 ;
        RECT 71.825 130.970 77.170 131.515 ;
        RECT 77.345 130.970 82.690 131.515 ;
        RECT 82.865 130.970 88.210 131.515 ;
        RECT 88.385 130.970 93.730 131.515 ;
        RECT 69.065 130.225 69.815 130.745 ;
        RECT 73.410 130.140 73.750 130.970 ;
        RECT 78.930 130.140 79.270 130.970 ;
        RECT 84.450 130.140 84.790 130.970 ;
        RECT 89.970 130.140 90.310 130.970 ;
        RECT 93.905 130.745 96.495 131.515 ;
        RECT 97.125 130.790 97.415 131.515 ;
        RECT 97.585 130.970 102.930 131.515 ;
        RECT 103.105 130.970 108.450 131.515 ;
        RECT 108.625 130.970 113.970 131.515 ;
        RECT 114.145 130.970 119.490 131.515 ;
        RECT 93.905 130.225 95.115 130.745 ;
        RECT 99.170 130.140 99.510 130.970 ;
        RECT 104.690 130.140 105.030 130.970 ;
        RECT 110.210 130.140 110.550 130.970 ;
        RECT 115.730 130.140 116.070 130.970 ;
        RECT 119.665 130.745 122.255 131.515 ;
        RECT 122.885 130.790 123.175 131.515 ;
        RECT 123.345 130.970 128.690 131.515 ;
        RECT 119.665 130.225 120.875 130.745 ;
        RECT 124.930 130.140 125.270 130.970 ;
        RECT 128.865 130.745 132.375 131.515 ;
        RECT 133.005 130.765 134.215 131.515 ;
        RECT 128.865 130.225 130.515 130.745 ;
        RECT 133.695 130.225 134.215 130.765 ;
        RECT 45.605 126.995 46.125 127.535 ;
        RECT 45.605 126.245 46.815 126.995 ;
        RECT 48.570 126.790 48.910 127.620 ;
        RECT 54.090 126.790 54.430 127.620 ;
        RECT 46.985 126.245 52.330 126.790 ;
        RECT 52.505 126.245 57.850 126.790 ;
        RECT 58.485 126.245 58.775 126.970 ;
        RECT 60.530 126.790 60.870 127.620 ;
        RECT 66.050 126.790 66.390 127.620 ;
        RECT 71.570 126.790 71.910 127.620 ;
        RECT 77.090 126.790 77.430 127.620 ;
        RECT 81.025 127.015 82.235 127.535 ;
        RECT 58.945 126.245 64.290 126.790 ;
        RECT 64.465 126.245 69.810 126.790 ;
        RECT 69.985 126.245 75.330 126.790 ;
        RECT 75.505 126.245 80.850 126.790 ;
        RECT 81.025 126.245 83.615 127.015 ;
        RECT 84.245 126.245 84.535 126.970 ;
        RECT 86.290 126.790 86.630 127.620 ;
        RECT 91.810 126.790 92.150 127.620 ;
        RECT 97.330 126.790 97.670 127.620 ;
        RECT 102.850 126.790 103.190 127.620 ;
        RECT 106.785 127.015 107.995 127.535 ;
        RECT 84.705 126.245 90.050 126.790 ;
        RECT 90.225 126.245 95.570 126.790 ;
        RECT 95.745 126.245 101.090 126.790 ;
        RECT 101.265 126.245 106.610 126.790 ;
        RECT 106.785 126.245 109.375 127.015 ;
        RECT 110.005 126.245 110.295 126.970 ;
        RECT 112.050 126.790 112.390 127.620 ;
        RECT 117.570 126.790 117.910 127.620 ;
        RECT 123.090 126.790 123.430 127.620 ;
        RECT 128.610 126.790 128.950 127.620 ;
        RECT 133.695 126.995 134.215 127.535 ;
        RECT 110.465 126.245 115.810 126.790 ;
        RECT 115.985 126.245 121.330 126.790 ;
        RECT 121.505 126.245 126.850 126.790 ;
        RECT 127.025 126.245 132.370 126.790 ;
        RECT 133.005 126.245 134.215 126.995 ;
        RECT 45.520 126.075 134.300 126.245 ;
        RECT 45.605 125.325 46.815 126.075 ;
        RECT 46.985 125.530 52.330 126.075 ;
        RECT 52.505 125.530 57.850 126.075 ;
        RECT 58.025 125.530 63.370 126.075 ;
        RECT 63.545 125.530 68.890 126.075 ;
        RECT 45.605 124.785 46.125 125.325 ;
        RECT 48.570 124.700 48.910 125.530 ;
        RECT 54.090 124.700 54.430 125.530 ;
        RECT 59.610 124.700 59.950 125.530 ;
        RECT 65.130 124.700 65.470 125.530 ;
        RECT 69.065 125.305 70.735 126.075 ;
        RECT 71.365 125.350 71.655 126.075 ;
        RECT 71.825 125.530 77.170 126.075 ;
        RECT 77.345 125.530 82.690 126.075 ;
        RECT 82.865 125.530 88.210 126.075 ;
        RECT 88.385 125.530 93.730 126.075 ;
        RECT 69.065 124.785 69.815 125.305 ;
        RECT 73.410 124.700 73.750 125.530 ;
        RECT 78.930 124.700 79.270 125.530 ;
        RECT 84.450 124.700 84.790 125.530 ;
        RECT 89.970 124.700 90.310 125.530 ;
        RECT 93.905 125.305 96.495 126.075 ;
        RECT 97.125 125.350 97.415 126.075 ;
        RECT 97.585 125.530 102.930 126.075 ;
        RECT 103.105 125.530 108.450 126.075 ;
        RECT 108.625 125.530 113.970 126.075 ;
        RECT 114.145 125.530 119.490 126.075 ;
        RECT 93.905 124.785 95.115 125.305 ;
        RECT 99.170 124.700 99.510 125.530 ;
        RECT 104.690 124.700 105.030 125.530 ;
        RECT 110.210 124.700 110.550 125.530 ;
        RECT 115.730 124.700 116.070 125.530 ;
        RECT 119.665 125.305 122.255 126.075 ;
        RECT 122.885 125.350 123.175 126.075 ;
        RECT 123.345 125.530 128.690 126.075 ;
        RECT 119.665 124.785 120.875 125.305 ;
        RECT 124.930 124.700 125.270 125.530 ;
        RECT 128.865 125.305 132.375 126.075 ;
        RECT 133.005 125.325 134.215 126.075 ;
        RECT 128.865 124.785 130.515 125.305 ;
        RECT 133.695 124.785 134.215 125.325 ;
        RECT 45.605 121.555 46.125 122.095 ;
        RECT 45.605 120.805 46.815 121.555 ;
        RECT 48.570 121.350 48.910 122.180 ;
        RECT 54.090 121.350 54.430 122.180 ;
        RECT 46.985 120.805 52.330 121.350 ;
        RECT 52.505 120.805 57.850 121.350 ;
        RECT 58.485 120.805 58.775 121.530 ;
        RECT 60.530 121.350 60.870 122.180 ;
        RECT 66.050 121.350 66.390 122.180 ;
        RECT 71.570 121.350 71.910 122.180 ;
        RECT 77.090 121.350 77.430 122.180 ;
        RECT 81.025 121.575 82.235 122.095 ;
        RECT 58.945 120.805 64.290 121.350 ;
        RECT 64.465 120.805 69.810 121.350 ;
        RECT 69.985 120.805 75.330 121.350 ;
        RECT 75.505 120.805 80.850 121.350 ;
        RECT 81.025 120.805 83.615 121.575 ;
        RECT 84.245 120.805 84.535 121.530 ;
        RECT 86.290 121.350 86.630 122.180 ;
        RECT 91.810 121.350 92.150 122.180 ;
        RECT 97.330 121.350 97.670 122.180 ;
        RECT 102.850 121.350 103.190 122.180 ;
        RECT 106.785 121.575 107.995 122.095 ;
        RECT 84.705 120.805 90.050 121.350 ;
        RECT 90.225 120.805 95.570 121.350 ;
        RECT 95.745 120.805 101.090 121.350 ;
        RECT 101.265 120.805 106.610 121.350 ;
        RECT 106.785 120.805 109.375 121.575 ;
        RECT 110.005 120.805 110.295 121.530 ;
        RECT 112.050 121.350 112.390 122.180 ;
        RECT 117.570 121.350 117.910 122.180 ;
        RECT 123.090 121.350 123.430 122.180 ;
        RECT 128.610 121.350 128.950 122.180 ;
        RECT 133.695 121.555 134.215 122.095 ;
        RECT 110.465 120.805 115.810 121.350 ;
        RECT 115.985 120.805 121.330 121.350 ;
        RECT 121.505 120.805 126.850 121.350 ;
        RECT 127.025 120.805 132.370 121.350 ;
        RECT 133.005 120.805 134.215 121.555 ;
        RECT 45.520 120.635 134.300 120.805 ;
        RECT 45.605 119.885 46.815 120.635 ;
        RECT 46.985 120.090 52.330 120.635 ;
        RECT 52.505 120.090 57.850 120.635 ;
        RECT 58.025 120.090 63.370 120.635 ;
        RECT 63.545 120.090 68.890 120.635 ;
        RECT 45.605 119.345 46.125 119.885 ;
        RECT 48.570 119.260 48.910 120.090 ;
        RECT 54.090 119.260 54.430 120.090 ;
        RECT 59.610 119.260 59.950 120.090 ;
        RECT 65.130 119.260 65.470 120.090 ;
        RECT 69.065 119.865 70.735 120.635 ;
        RECT 71.365 119.910 71.655 120.635 ;
        RECT 71.825 120.090 77.170 120.635 ;
        RECT 77.345 120.090 82.690 120.635 ;
        RECT 82.865 120.090 88.210 120.635 ;
        RECT 88.385 120.090 93.730 120.635 ;
        RECT 69.065 119.345 69.815 119.865 ;
        RECT 73.410 119.260 73.750 120.090 ;
        RECT 78.930 119.260 79.270 120.090 ;
        RECT 84.450 119.260 84.790 120.090 ;
        RECT 89.970 119.260 90.310 120.090 ;
        RECT 93.905 119.865 96.495 120.635 ;
        RECT 97.125 119.910 97.415 120.635 ;
        RECT 97.585 120.090 102.930 120.635 ;
        RECT 103.105 120.090 108.450 120.635 ;
        RECT 108.625 120.090 113.970 120.635 ;
        RECT 114.145 120.090 119.490 120.635 ;
        RECT 93.905 119.345 95.115 119.865 ;
        RECT 99.170 119.260 99.510 120.090 ;
        RECT 104.690 119.260 105.030 120.090 ;
        RECT 110.210 119.260 110.550 120.090 ;
        RECT 115.730 119.260 116.070 120.090 ;
        RECT 119.665 119.865 122.255 120.635 ;
        RECT 122.885 119.910 123.175 120.635 ;
        RECT 123.345 120.090 128.690 120.635 ;
        RECT 119.665 119.345 120.875 119.865 ;
        RECT 124.930 119.260 125.270 120.090 ;
        RECT 128.865 119.865 132.375 120.635 ;
        RECT 133.005 119.885 134.215 120.635 ;
        RECT 128.865 119.345 130.515 119.865 ;
        RECT 133.695 119.345 134.215 119.885 ;
        RECT 45.605 116.115 46.125 116.655 ;
        RECT 45.605 115.365 46.815 116.115 ;
        RECT 48.570 115.910 48.910 116.740 ;
        RECT 54.090 115.910 54.430 116.740 ;
        RECT 46.985 115.365 52.330 115.910 ;
        RECT 52.505 115.365 57.850 115.910 ;
        RECT 58.485 115.365 58.775 116.090 ;
        RECT 60.530 115.910 60.870 116.740 ;
        RECT 66.050 115.910 66.390 116.740 ;
        RECT 71.570 115.910 71.910 116.740 ;
        RECT 77.090 115.910 77.430 116.740 ;
        RECT 81.025 116.135 82.235 116.655 ;
        RECT 58.945 115.365 64.290 115.910 ;
        RECT 64.465 115.365 69.810 115.910 ;
        RECT 69.985 115.365 75.330 115.910 ;
        RECT 75.505 115.365 80.850 115.910 ;
        RECT 81.025 115.365 83.615 116.135 ;
        RECT 84.245 115.365 84.535 116.090 ;
        RECT 86.290 115.910 86.630 116.740 ;
        RECT 91.810 115.910 92.150 116.740 ;
        RECT 97.330 115.910 97.670 116.740 ;
        RECT 102.850 115.910 103.190 116.740 ;
        RECT 106.785 116.135 107.995 116.655 ;
        RECT 84.705 115.365 90.050 115.910 ;
        RECT 90.225 115.365 95.570 115.910 ;
        RECT 95.745 115.365 101.090 115.910 ;
        RECT 101.265 115.365 106.610 115.910 ;
        RECT 106.785 115.365 109.375 116.135 ;
        RECT 110.005 115.365 110.295 116.090 ;
        RECT 112.050 115.910 112.390 116.740 ;
        RECT 117.570 115.910 117.910 116.740 ;
        RECT 123.090 115.910 123.430 116.740 ;
        RECT 128.610 115.910 128.950 116.740 ;
        RECT 133.695 116.115 134.215 116.655 ;
        RECT 110.465 115.365 115.810 115.910 ;
        RECT 115.985 115.365 121.330 115.910 ;
        RECT 121.505 115.365 126.850 115.910 ;
        RECT 127.025 115.365 132.370 115.910 ;
        RECT 133.005 115.365 134.215 116.115 ;
        RECT 45.520 115.195 134.300 115.365 ;
        RECT 45.605 114.445 46.815 115.195 ;
        RECT 46.985 114.650 52.330 115.195 ;
        RECT 52.505 114.650 57.850 115.195 ;
        RECT 58.025 114.650 63.370 115.195 ;
        RECT 63.545 114.650 68.890 115.195 ;
        RECT 45.605 113.905 46.125 114.445 ;
        RECT 48.570 113.820 48.910 114.650 ;
        RECT 54.090 113.820 54.430 114.650 ;
        RECT 59.610 113.820 59.950 114.650 ;
        RECT 65.130 113.820 65.470 114.650 ;
        RECT 69.065 114.425 70.735 115.195 ;
        RECT 71.365 114.470 71.655 115.195 ;
        RECT 71.825 114.650 77.170 115.195 ;
        RECT 77.345 114.650 82.690 115.195 ;
        RECT 82.865 114.650 88.210 115.195 ;
        RECT 88.385 114.650 93.730 115.195 ;
        RECT 69.065 113.905 69.815 114.425 ;
        RECT 73.410 113.820 73.750 114.650 ;
        RECT 78.930 113.820 79.270 114.650 ;
        RECT 84.450 113.820 84.790 114.650 ;
        RECT 89.970 113.820 90.310 114.650 ;
        RECT 93.905 114.425 96.495 115.195 ;
        RECT 97.125 114.470 97.415 115.195 ;
        RECT 97.585 114.650 102.930 115.195 ;
        RECT 103.105 114.650 108.450 115.195 ;
        RECT 108.625 114.650 113.970 115.195 ;
        RECT 114.145 114.650 119.490 115.195 ;
        RECT 93.905 113.905 95.115 114.425 ;
        RECT 99.170 113.820 99.510 114.650 ;
        RECT 104.690 113.820 105.030 114.650 ;
        RECT 110.210 113.820 110.550 114.650 ;
        RECT 115.730 113.820 116.070 114.650 ;
        RECT 119.665 114.425 122.255 115.195 ;
        RECT 122.885 114.470 123.175 115.195 ;
        RECT 123.345 114.650 128.690 115.195 ;
        RECT 119.665 113.905 120.875 114.425 ;
        RECT 124.930 113.820 125.270 114.650 ;
        RECT 128.865 114.425 132.375 115.195 ;
        RECT 133.005 114.445 134.215 115.195 ;
        RECT 128.865 113.905 130.515 114.425 ;
        RECT 133.695 113.905 134.215 114.445 ;
        RECT 45.605 110.675 46.125 111.215 ;
        RECT 45.605 109.925 46.815 110.675 ;
        RECT 48.570 110.470 48.910 111.300 ;
        RECT 54.090 110.470 54.430 111.300 ;
        RECT 46.985 109.925 52.330 110.470 ;
        RECT 52.505 109.925 57.850 110.470 ;
        RECT 58.485 109.925 58.775 110.650 ;
        RECT 60.530 110.470 60.870 111.300 ;
        RECT 66.050 110.470 66.390 111.300 ;
        RECT 71.570 110.470 71.910 111.300 ;
        RECT 77.090 110.470 77.430 111.300 ;
        RECT 81.025 110.695 82.235 111.215 ;
        RECT 58.945 109.925 64.290 110.470 ;
        RECT 64.465 109.925 69.810 110.470 ;
        RECT 69.985 109.925 75.330 110.470 ;
        RECT 75.505 109.925 80.850 110.470 ;
        RECT 81.025 109.925 83.615 110.695 ;
        RECT 84.245 109.925 84.535 110.650 ;
        RECT 86.290 110.470 86.630 111.300 ;
        RECT 91.810 110.470 92.150 111.300 ;
        RECT 97.330 110.470 97.670 111.300 ;
        RECT 102.850 110.470 103.190 111.300 ;
        RECT 106.785 110.695 107.995 111.215 ;
        RECT 84.705 109.925 90.050 110.470 ;
        RECT 90.225 109.925 95.570 110.470 ;
        RECT 95.745 109.925 101.090 110.470 ;
        RECT 101.265 109.925 106.610 110.470 ;
        RECT 106.785 109.925 109.375 110.695 ;
        RECT 110.005 109.925 110.295 110.650 ;
        RECT 112.050 110.470 112.390 111.300 ;
        RECT 117.570 110.470 117.910 111.300 ;
        RECT 123.090 110.470 123.430 111.300 ;
        RECT 128.610 110.470 128.950 111.300 ;
        RECT 133.695 110.675 134.215 111.215 ;
        RECT 110.465 109.925 115.810 110.470 ;
        RECT 115.985 109.925 121.330 110.470 ;
        RECT 121.505 109.925 126.850 110.470 ;
        RECT 127.025 109.925 132.370 110.470 ;
        RECT 133.005 109.925 134.215 110.675 ;
        RECT 45.520 109.755 134.300 109.925 ;
        RECT 45.605 109.005 46.815 109.755 ;
        RECT 46.985 109.210 52.330 109.755 ;
        RECT 52.505 109.210 57.850 109.755 ;
        RECT 45.605 108.465 46.125 109.005 ;
        RECT 48.570 108.380 48.910 109.210 ;
        RECT 54.090 108.380 54.430 109.210 ;
        RECT 58.025 108.985 59.695 109.755 ;
        RECT 58.025 108.465 58.775 108.985 ;
        RECT 60.365 108.935 60.595 109.755 ;
        RECT 61.265 108.935 61.475 109.755 ;
        RECT 62.180 109.375 62.510 109.755 ;
        RECT 63.110 108.915 63.370 109.755 ;
        RECT 63.545 109.210 68.890 109.755 ;
        RECT 65.130 108.380 65.470 109.210 ;
        RECT 69.065 108.985 70.735 109.755 ;
        RECT 71.365 109.030 71.655 109.755 ;
        RECT 71.825 109.210 77.170 109.755 ;
        RECT 77.345 109.210 82.690 109.755 ;
        RECT 82.865 109.210 88.210 109.755 ;
        RECT 88.385 109.210 93.730 109.755 ;
        RECT 69.065 108.465 69.815 108.985 ;
        RECT 73.410 108.380 73.750 109.210 ;
        RECT 78.930 108.380 79.270 109.210 ;
        RECT 84.450 108.380 84.790 109.210 ;
        RECT 89.970 108.380 90.310 109.210 ;
        RECT 93.905 108.985 96.495 109.755 ;
        RECT 97.125 109.030 97.415 109.755 ;
        RECT 97.585 109.210 102.930 109.755 ;
        RECT 103.105 109.210 108.450 109.755 ;
        RECT 108.625 109.210 113.970 109.755 ;
        RECT 114.145 109.210 119.490 109.755 ;
        RECT 93.905 108.465 95.115 108.985 ;
        RECT 99.170 108.380 99.510 109.210 ;
        RECT 104.690 108.380 105.030 109.210 ;
        RECT 110.210 108.380 110.550 109.210 ;
        RECT 115.730 108.380 116.070 109.210 ;
        RECT 119.665 108.985 122.255 109.755 ;
        RECT 122.885 109.030 123.175 109.755 ;
        RECT 123.345 109.210 128.690 109.755 ;
        RECT 119.665 108.465 120.875 108.985 ;
        RECT 124.930 108.380 125.270 109.210 ;
        RECT 128.865 108.985 132.375 109.755 ;
        RECT 133.005 109.005 134.215 109.755 ;
        RECT 128.865 108.465 130.515 108.985 ;
        RECT 133.695 108.465 134.215 109.005 ;
        RECT 45.605 105.235 46.125 105.775 ;
        RECT 46.985 105.255 48.635 105.775 ;
        RECT 45.605 104.485 46.815 105.235 ;
        RECT 46.985 104.485 50.495 105.255 ;
        RECT 51.185 104.485 51.395 105.305 ;
        RECT 52.065 104.485 52.295 105.305 ;
        RECT 52.505 104.485 52.815 105.285 ;
        RECT 54.525 104.485 55.285 104.965 ;
        RECT 56.635 104.485 56.965 104.845 ;
        RECT 58.485 104.485 58.775 105.210 ;
        RECT 60.530 105.030 60.870 105.860 ;
        RECT 66.050 105.030 66.390 105.860 ;
        RECT 71.570 105.030 71.910 105.860 ;
        RECT 77.090 105.030 77.430 105.860 ;
        RECT 81.025 105.255 82.235 105.775 ;
        RECT 58.945 104.485 64.290 105.030 ;
        RECT 64.465 104.485 69.810 105.030 ;
        RECT 69.985 104.485 75.330 105.030 ;
        RECT 75.505 104.485 80.850 105.030 ;
        RECT 81.025 104.485 83.615 105.255 ;
        RECT 84.245 104.485 84.535 105.210 ;
        RECT 86.290 105.030 86.630 105.860 ;
        RECT 91.810 105.030 92.150 105.860 ;
        RECT 97.330 105.030 97.670 105.860 ;
        RECT 102.850 105.030 103.190 105.860 ;
        RECT 106.785 105.255 107.995 105.775 ;
        RECT 84.705 104.485 90.050 105.030 ;
        RECT 90.225 104.485 95.570 105.030 ;
        RECT 95.745 104.485 101.090 105.030 ;
        RECT 101.265 104.485 106.610 105.030 ;
        RECT 106.785 104.485 109.375 105.255 ;
        RECT 110.005 104.485 110.295 105.210 ;
        RECT 112.050 105.030 112.390 105.860 ;
        RECT 117.570 105.030 117.910 105.860 ;
        RECT 123.090 105.030 123.430 105.860 ;
        RECT 128.610 105.030 128.950 105.860 ;
        RECT 133.695 105.235 134.215 105.775 ;
        RECT 110.465 104.485 115.810 105.030 ;
        RECT 115.985 104.485 121.330 105.030 ;
        RECT 121.505 104.485 126.850 105.030 ;
        RECT 127.025 104.485 132.370 105.030 ;
        RECT 133.005 104.485 134.215 105.235 ;
        RECT 45.520 104.315 134.300 104.485 ;
        RECT 45.605 103.565 46.815 104.315 ;
        RECT 47.425 103.935 47.755 104.315 ;
        RECT 48.365 103.770 53.710 104.315 ;
        RECT 55.315 103.855 55.485 104.315 ;
        RECT 57.535 103.805 57.870 104.315 ;
        RECT 59.360 103.915 59.690 104.315 ;
        RECT 61.245 103.770 66.590 104.315 ;
        RECT 45.605 103.025 46.125 103.565 ;
        RECT 49.950 102.940 50.290 103.770 ;
        RECT 62.830 102.940 63.170 103.770 ;
        RECT 66.765 103.545 70.275 104.315 ;
        RECT 71.365 103.590 71.655 104.315 ;
        RECT 71.825 103.770 77.170 104.315 ;
        RECT 77.345 103.770 82.690 104.315 ;
        RECT 82.865 103.770 88.210 104.315 ;
        RECT 88.385 103.770 93.730 104.315 ;
        RECT 66.765 103.025 68.415 103.545 ;
        RECT 73.410 102.940 73.750 103.770 ;
        RECT 78.930 102.940 79.270 103.770 ;
        RECT 84.450 102.940 84.790 103.770 ;
        RECT 89.970 102.940 90.310 103.770 ;
        RECT 93.905 103.545 96.495 104.315 ;
        RECT 97.125 103.590 97.415 104.315 ;
        RECT 97.585 103.770 102.930 104.315 ;
        RECT 103.105 103.770 108.450 104.315 ;
        RECT 108.625 103.770 113.970 104.315 ;
        RECT 114.145 103.770 119.490 104.315 ;
        RECT 93.905 103.025 95.115 103.545 ;
        RECT 99.170 102.940 99.510 103.770 ;
        RECT 104.690 102.940 105.030 103.770 ;
        RECT 110.210 102.940 110.550 103.770 ;
        RECT 115.730 102.940 116.070 103.770 ;
        RECT 119.665 103.545 122.255 104.315 ;
        RECT 122.885 103.590 123.175 104.315 ;
        RECT 123.345 103.770 128.690 104.315 ;
        RECT 119.665 103.025 120.875 103.545 ;
        RECT 124.930 102.940 125.270 103.770 ;
        RECT 128.865 103.545 132.375 104.315 ;
        RECT 133.005 103.565 134.215 104.315 ;
        RECT 128.865 103.025 130.515 103.545 ;
        RECT 133.695 103.025 134.215 103.565 ;
        RECT 45.605 99.795 46.125 100.335 ;
        RECT 45.605 99.045 46.815 99.795 ;
        RECT 49.950 99.590 50.290 100.420 ;
        RECT 53.885 99.815 55.535 100.335 ;
        RECT 47.425 99.045 47.755 99.425 ;
        RECT 48.365 99.045 53.710 99.590 ;
        RECT 53.885 99.045 57.395 99.815 ;
        RECT 58.485 99.045 58.775 99.770 ;
        RECT 60.530 99.590 60.870 100.420 ;
        RECT 66.050 99.590 66.390 100.420 ;
        RECT 71.570 99.590 71.910 100.420 ;
        RECT 77.090 99.590 77.430 100.420 ;
        RECT 81.025 99.815 82.235 100.335 ;
        RECT 58.945 99.045 64.290 99.590 ;
        RECT 64.465 99.045 69.810 99.590 ;
        RECT 69.985 99.045 75.330 99.590 ;
        RECT 75.505 99.045 80.850 99.590 ;
        RECT 81.025 99.045 83.615 99.815 ;
        RECT 84.245 99.045 84.535 99.770 ;
        RECT 86.290 99.590 86.630 100.420 ;
        RECT 91.810 99.590 92.150 100.420 ;
        RECT 97.330 99.590 97.670 100.420 ;
        RECT 102.850 99.590 103.190 100.420 ;
        RECT 106.785 99.815 107.995 100.335 ;
        RECT 84.705 99.045 90.050 99.590 ;
        RECT 90.225 99.045 95.570 99.590 ;
        RECT 95.745 99.045 101.090 99.590 ;
        RECT 101.265 99.045 106.610 99.590 ;
        RECT 106.785 99.045 109.375 99.815 ;
        RECT 110.005 99.045 110.295 99.770 ;
        RECT 112.050 99.590 112.390 100.420 ;
        RECT 117.570 99.590 117.910 100.420 ;
        RECT 123.090 99.590 123.430 100.420 ;
        RECT 128.610 99.590 128.950 100.420 ;
        RECT 133.695 99.795 134.215 100.335 ;
        RECT 110.465 99.045 115.810 99.590 ;
        RECT 115.985 99.045 121.330 99.590 ;
        RECT 121.505 99.045 126.850 99.590 ;
        RECT 127.025 99.045 132.370 99.590 ;
        RECT 133.005 99.045 134.215 99.795 ;
        RECT 45.520 98.875 134.300 99.045 ;
        RECT 45.605 98.125 46.815 98.875 ;
        RECT 46.985 98.330 52.330 98.875 ;
        RECT 45.605 97.585 46.125 98.125 ;
        RECT 48.570 97.500 48.910 98.330 ;
        RECT 52.505 98.105 55.095 98.875 ;
        RECT 56.165 98.495 56.495 98.875 ;
        RECT 57.105 98.330 62.450 98.875 ;
        RECT 62.625 98.330 67.970 98.875 ;
        RECT 52.505 97.585 53.715 98.105 ;
        RECT 58.690 97.500 59.030 98.330 ;
        RECT 64.210 97.500 64.550 98.330 ;
        RECT 68.145 98.105 70.735 98.875 ;
        RECT 71.365 98.150 71.655 98.875 ;
        RECT 71.825 98.330 77.170 98.875 ;
        RECT 77.345 98.330 82.690 98.875 ;
        RECT 82.865 98.330 88.210 98.875 ;
        RECT 88.385 98.330 93.730 98.875 ;
        RECT 68.145 97.585 69.355 98.105 ;
        RECT 73.410 97.500 73.750 98.330 ;
        RECT 78.930 97.500 79.270 98.330 ;
        RECT 84.450 97.500 84.790 98.330 ;
        RECT 89.970 97.500 90.310 98.330 ;
        RECT 93.905 98.105 96.495 98.875 ;
        RECT 97.125 98.150 97.415 98.875 ;
        RECT 97.585 98.330 102.930 98.875 ;
        RECT 103.105 98.330 108.450 98.875 ;
        RECT 108.625 98.330 113.970 98.875 ;
        RECT 114.145 98.330 119.490 98.875 ;
        RECT 93.905 97.585 95.115 98.105 ;
        RECT 99.170 97.500 99.510 98.330 ;
        RECT 104.690 97.500 105.030 98.330 ;
        RECT 110.210 97.500 110.550 98.330 ;
        RECT 115.730 97.500 116.070 98.330 ;
        RECT 119.665 98.105 122.255 98.875 ;
        RECT 122.885 98.150 123.175 98.875 ;
        RECT 123.345 98.330 128.690 98.875 ;
        RECT 119.665 97.585 120.875 98.105 ;
        RECT 124.930 97.500 125.270 98.330 ;
        RECT 128.865 98.105 132.375 98.875 ;
        RECT 133.005 98.125 134.215 98.875 ;
        RECT 128.865 97.585 130.515 98.105 ;
        RECT 133.695 97.585 134.215 98.125 ;
        RECT 45.605 94.355 46.125 94.895 ;
        RECT 45.605 93.605 46.815 94.355 ;
        RECT 48.570 94.150 48.910 94.980 ;
        RECT 52.505 94.375 54.155 94.895 ;
        RECT 46.985 93.605 52.330 94.150 ;
        RECT 52.505 93.605 56.015 94.375 ;
        RECT 57.545 93.605 57.855 94.405 ;
        RECT 58.485 93.605 58.775 94.330 ;
        RECT 60.530 94.150 60.870 94.980 ;
        RECT 66.050 94.150 66.390 94.980 ;
        RECT 71.570 94.150 71.910 94.980 ;
        RECT 77.090 94.150 77.430 94.980 ;
        RECT 81.025 94.375 82.235 94.895 ;
        RECT 58.945 93.605 64.290 94.150 ;
        RECT 64.465 93.605 69.810 94.150 ;
        RECT 69.985 93.605 75.330 94.150 ;
        RECT 75.505 93.605 80.850 94.150 ;
        RECT 81.025 93.605 83.615 94.375 ;
        RECT 84.245 93.605 84.535 94.330 ;
        RECT 86.290 94.150 86.630 94.980 ;
        RECT 91.810 94.150 92.150 94.980 ;
        RECT 97.330 94.150 97.670 94.980 ;
        RECT 102.850 94.150 103.190 94.980 ;
        RECT 106.785 94.375 107.995 94.895 ;
        RECT 84.705 93.605 90.050 94.150 ;
        RECT 90.225 93.605 95.570 94.150 ;
        RECT 95.745 93.605 101.090 94.150 ;
        RECT 101.265 93.605 106.610 94.150 ;
        RECT 106.785 93.605 109.375 94.375 ;
        RECT 110.005 93.605 110.295 94.330 ;
        RECT 112.050 94.150 112.390 94.980 ;
        RECT 117.570 94.150 117.910 94.980 ;
        RECT 123.090 94.150 123.430 94.980 ;
        RECT 128.610 94.150 128.950 94.980 ;
        RECT 133.695 94.355 134.215 94.895 ;
        RECT 110.465 93.605 115.810 94.150 ;
        RECT 115.985 93.605 121.330 94.150 ;
        RECT 121.505 93.605 126.850 94.150 ;
        RECT 127.025 93.605 132.370 94.150 ;
        RECT 133.005 93.605 134.215 94.355 ;
        RECT 45.520 93.435 134.300 93.605 ;
        RECT 45.605 92.685 46.815 93.435 ;
        RECT 45.605 92.145 46.125 92.685 ;
        RECT 46.985 92.665 50.495 93.435 ;
        RECT 52.325 92.900 52.835 93.435 ;
        RECT 54.795 93.035 55.125 93.435 ;
        RECT 56.155 93.035 56.485 93.435 ;
        RECT 58.445 92.900 58.955 93.435 ;
        RECT 46.985 92.145 48.635 92.665 ;
        RECT 59.905 92.615 60.135 93.435 ;
        RECT 60.805 92.615 61.015 93.435 ;
        RECT 61.285 92.615 61.515 93.435 ;
        RECT 62.185 92.615 62.395 93.435 ;
        RECT 62.625 92.890 67.970 93.435 ;
        RECT 64.210 92.060 64.550 92.890 ;
        RECT 68.145 92.665 70.735 93.435 ;
        RECT 71.365 92.710 71.655 93.435 ;
        RECT 71.825 92.890 77.170 93.435 ;
        RECT 77.345 92.890 82.690 93.435 ;
        RECT 82.865 92.890 88.210 93.435 ;
        RECT 88.385 92.890 93.730 93.435 ;
        RECT 68.145 92.145 69.355 92.665 ;
        RECT 73.410 92.060 73.750 92.890 ;
        RECT 78.930 92.060 79.270 92.890 ;
        RECT 84.450 92.060 84.790 92.890 ;
        RECT 89.970 92.060 90.310 92.890 ;
        RECT 93.905 92.665 96.495 93.435 ;
        RECT 97.125 92.710 97.415 93.435 ;
        RECT 97.585 92.890 102.930 93.435 ;
        RECT 103.105 92.890 108.450 93.435 ;
        RECT 108.625 92.890 113.970 93.435 ;
        RECT 114.145 92.890 119.490 93.435 ;
        RECT 93.905 92.145 95.115 92.665 ;
        RECT 99.170 92.060 99.510 92.890 ;
        RECT 104.690 92.060 105.030 92.890 ;
        RECT 110.210 92.060 110.550 92.890 ;
        RECT 115.730 92.060 116.070 92.890 ;
        RECT 119.665 92.665 122.255 93.435 ;
        RECT 122.885 92.710 123.175 93.435 ;
        RECT 123.345 92.890 128.690 93.435 ;
        RECT 119.665 92.145 120.875 92.665 ;
        RECT 124.930 92.060 125.270 92.890 ;
        RECT 128.865 92.665 132.375 93.435 ;
        RECT 133.005 92.685 134.215 93.435 ;
        RECT 128.865 92.145 130.515 92.665 ;
        RECT 133.695 92.145 134.215 92.685 ;
        RECT 45.605 88.915 46.125 89.455 ;
        RECT 45.605 88.165 46.815 88.915 ;
        RECT 48.570 88.710 48.910 89.540 ;
        RECT 52.505 88.935 53.715 89.455 ;
        RECT 46.985 88.165 52.330 88.710 ;
        RECT 52.505 88.165 55.095 88.935 ;
        RECT 55.705 88.165 56.035 88.545 ;
        RECT 56.685 88.165 56.915 88.985 ;
        RECT 57.585 88.165 57.795 88.985 ;
        RECT 58.485 88.165 58.775 88.890 ;
        RECT 60.530 88.710 60.870 89.540 ;
        RECT 66.050 88.710 66.390 89.540 ;
        RECT 71.570 88.710 71.910 89.540 ;
        RECT 77.090 88.710 77.430 89.540 ;
        RECT 81.025 88.935 82.235 89.455 ;
        RECT 58.945 88.165 64.290 88.710 ;
        RECT 64.465 88.165 69.810 88.710 ;
        RECT 69.985 88.165 75.330 88.710 ;
        RECT 75.505 88.165 80.850 88.710 ;
        RECT 81.025 88.165 83.615 88.935 ;
        RECT 84.245 88.165 84.535 88.890 ;
        RECT 86.290 88.710 86.630 89.540 ;
        RECT 91.810 88.710 92.150 89.540 ;
        RECT 97.330 88.710 97.670 89.540 ;
        RECT 102.850 88.710 103.190 89.540 ;
        RECT 106.785 88.935 107.995 89.455 ;
        RECT 84.705 88.165 90.050 88.710 ;
        RECT 90.225 88.165 95.570 88.710 ;
        RECT 95.745 88.165 101.090 88.710 ;
        RECT 101.265 88.165 106.610 88.710 ;
        RECT 106.785 88.165 109.375 88.935 ;
        RECT 110.005 88.165 110.295 88.890 ;
        RECT 112.050 88.710 112.390 89.540 ;
        RECT 117.570 88.710 117.910 89.540 ;
        RECT 123.090 88.710 123.430 89.540 ;
        RECT 128.610 88.710 128.950 89.540 ;
        RECT 133.695 88.915 134.215 89.455 ;
        RECT 110.465 88.165 115.810 88.710 ;
        RECT 115.985 88.165 121.330 88.710 ;
        RECT 121.505 88.165 126.850 88.710 ;
        RECT 127.025 88.165 132.370 88.710 ;
        RECT 133.005 88.165 134.215 88.915 ;
        RECT 45.520 87.995 134.300 88.165 ;
        RECT 45.605 87.245 46.815 87.995 ;
        RECT 46.985 87.450 52.330 87.995 ;
        RECT 52.505 87.450 57.850 87.995 ;
        RECT 58.025 87.450 63.370 87.995 ;
        RECT 63.545 87.450 68.890 87.995 ;
        RECT 45.605 86.705 46.125 87.245 ;
        RECT 48.570 86.620 48.910 87.450 ;
        RECT 54.090 86.620 54.430 87.450 ;
        RECT 59.610 86.620 59.950 87.450 ;
        RECT 65.130 86.620 65.470 87.450 ;
        RECT 69.065 87.225 70.735 87.995 ;
        RECT 71.365 87.270 71.655 87.995 ;
        RECT 71.825 87.450 77.170 87.995 ;
        RECT 77.345 87.450 82.690 87.995 ;
        RECT 82.865 87.450 88.210 87.995 ;
        RECT 88.385 87.450 93.730 87.995 ;
        RECT 69.065 86.705 69.815 87.225 ;
        RECT 73.410 86.620 73.750 87.450 ;
        RECT 78.930 86.620 79.270 87.450 ;
        RECT 84.450 86.620 84.790 87.450 ;
        RECT 89.970 86.620 90.310 87.450 ;
        RECT 93.905 87.225 96.495 87.995 ;
        RECT 97.125 87.270 97.415 87.995 ;
        RECT 97.585 87.450 102.930 87.995 ;
        RECT 103.105 87.450 108.450 87.995 ;
        RECT 108.625 87.450 113.970 87.995 ;
        RECT 114.145 87.450 119.490 87.995 ;
        RECT 93.905 86.705 95.115 87.225 ;
        RECT 99.170 86.620 99.510 87.450 ;
        RECT 104.690 86.620 105.030 87.450 ;
        RECT 110.210 86.620 110.550 87.450 ;
        RECT 115.730 86.620 116.070 87.450 ;
        RECT 119.665 87.225 122.255 87.995 ;
        RECT 122.885 87.270 123.175 87.995 ;
        RECT 123.345 87.450 128.690 87.995 ;
        RECT 119.665 86.705 120.875 87.225 ;
        RECT 124.930 86.620 125.270 87.450 ;
        RECT 128.865 87.225 132.375 87.995 ;
        RECT 133.005 87.245 134.215 87.995 ;
        RECT 128.865 86.705 130.515 87.225 ;
        RECT 133.695 86.705 134.215 87.245 ;
        RECT 45.605 83.475 46.125 84.015 ;
        RECT 45.605 82.725 46.815 83.475 ;
        RECT 48.570 83.270 48.910 84.100 ;
        RECT 54.090 83.270 54.430 84.100 ;
        RECT 46.985 82.725 52.330 83.270 ;
        RECT 52.505 82.725 57.850 83.270 ;
        RECT 58.485 82.725 58.775 83.450 ;
        RECT 60.530 83.270 60.870 84.100 ;
        RECT 66.050 83.270 66.390 84.100 ;
        RECT 71.570 83.270 71.910 84.100 ;
        RECT 77.090 83.270 77.430 84.100 ;
        RECT 81.025 83.495 82.235 84.015 ;
        RECT 58.945 82.725 64.290 83.270 ;
        RECT 64.465 82.725 69.810 83.270 ;
        RECT 69.985 82.725 75.330 83.270 ;
        RECT 75.505 82.725 80.850 83.270 ;
        RECT 81.025 82.725 83.615 83.495 ;
        RECT 84.245 82.725 84.535 83.450 ;
        RECT 86.290 83.270 86.630 84.100 ;
        RECT 91.810 83.270 92.150 84.100 ;
        RECT 97.330 83.270 97.670 84.100 ;
        RECT 102.850 83.270 103.190 84.100 ;
        RECT 106.785 83.495 107.995 84.015 ;
        RECT 84.705 82.725 90.050 83.270 ;
        RECT 90.225 82.725 95.570 83.270 ;
        RECT 95.745 82.725 101.090 83.270 ;
        RECT 101.265 82.725 106.610 83.270 ;
        RECT 106.785 82.725 109.375 83.495 ;
        RECT 110.005 82.725 110.295 83.450 ;
        RECT 112.050 83.270 112.390 84.100 ;
        RECT 117.570 83.270 117.910 84.100 ;
        RECT 123.090 83.270 123.430 84.100 ;
        RECT 128.610 83.270 128.950 84.100 ;
        RECT 133.695 83.475 134.215 84.015 ;
        RECT 110.465 82.725 115.810 83.270 ;
        RECT 115.985 82.725 121.330 83.270 ;
        RECT 121.505 82.725 126.850 83.270 ;
        RECT 127.025 82.725 132.370 83.270 ;
        RECT 133.005 82.725 134.215 83.475 ;
        RECT 45.520 82.555 134.300 82.725 ;
        RECT 45.605 81.805 46.815 82.555 ;
        RECT 46.985 82.010 52.330 82.555 ;
        RECT 52.505 82.010 57.850 82.555 ;
        RECT 58.025 82.010 63.370 82.555 ;
        RECT 63.545 82.010 68.890 82.555 ;
        RECT 45.605 81.265 46.125 81.805 ;
        RECT 48.570 81.180 48.910 82.010 ;
        RECT 54.090 81.180 54.430 82.010 ;
        RECT 59.610 81.180 59.950 82.010 ;
        RECT 65.130 81.180 65.470 82.010 ;
        RECT 69.065 81.785 70.735 82.555 ;
        RECT 71.365 81.830 71.655 82.555 ;
        RECT 71.825 82.010 77.170 82.555 ;
        RECT 77.345 82.010 82.690 82.555 ;
        RECT 82.865 82.010 88.210 82.555 ;
        RECT 88.385 82.010 93.730 82.555 ;
        RECT 69.065 81.265 69.815 81.785 ;
        RECT 73.410 81.180 73.750 82.010 ;
        RECT 78.930 81.180 79.270 82.010 ;
        RECT 84.450 81.180 84.790 82.010 ;
        RECT 89.970 81.180 90.310 82.010 ;
        RECT 93.905 81.785 96.495 82.555 ;
        RECT 97.125 81.830 97.415 82.555 ;
        RECT 97.585 82.010 102.930 82.555 ;
        RECT 103.105 82.010 108.450 82.555 ;
        RECT 108.625 82.010 113.970 82.555 ;
        RECT 114.145 82.010 119.490 82.555 ;
        RECT 93.905 81.265 95.115 81.785 ;
        RECT 99.170 81.180 99.510 82.010 ;
        RECT 104.690 81.180 105.030 82.010 ;
        RECT 110.210 81.180 110.550 82.010 ;
        RECT 115.730 81.180 116.070 82.010 ;
        RECT 119.665 81.785 122.255 82.555 ;
        RECT 122.885 81.830 123.175 82.555 ;
        RECT 123.345 82.010 128.690 82.555 ;
        RECT 119.665 81.265 120.875 81.785 ;
        RECT 124.930 81.180 125.270 82.010 ;
        RECT 128.865 81.785 132.375 82.555 ;
        RECT 133.005 81.805 134.215 82.555 ;
        RECT 128.865 81.265 130.515 81.785 ;
        RECT 133.695 81.265 134.215 81.805 ;
        RECT 45.605 78.035 46.125 78.575 ;
        RECT 45.605 77.285 46.815 78.035 ;
        RECT 48.570 77.830 48.910 78.660 ;
        RECT 54.090 77.830 54.430 78.660 ;
        RECT 46.985 77.285 52.330 77.830 ;
        RECT 52.505 77.285 57.850 77.830 ;
        RECT 58.485 77.285 58.775 78.010 ;
        RECT 60.530 77.830 60.870 78.660 ;
        RECT 66.050 77.830 66.390 78.660 ;
        RECT 71.570 77.830 71.910 78.660 ;
        RECT 77.090 77.830 77.430 78.660 ;
        RECT 81.025 78.055 82.235 78.575 ;
        RECT 58.945 77.285 64.290 77.830 ;
        RECT 64.465 77.285 69.810 77.830 ;
        RECT 69.985 77.285 75.330 77.830 ;
        RECT 75.505 77.285 80.850 77.830 ;
        RECT 81.025 77.285 83.615 78.055 ;
        RECT 84.245 77.285 84.535 78.010 ;
        RECT 86.290 77.830 86.630 78.660 ;
        RECT 91.810 77.830 92.150 78.660 ;
        RECT 97.330 77.830 97.670 78.660 ;
        RECT 102.850 77.830 103.190 78.660 ;
        RECT 106.785 78.055 107.995 78.575 ;
        RECT 84.705 77.285 90.050 77.830 ;
        RECT 90.225 77.285 95.570 77.830 ;
        RECT 95.745 77.285 101.090 77.830 ;
        RECT 101.265 77.285 106.610 77.830 ;
        RECT 106.785 77.285 109.375 78.055 ;
        RECT 110.005 77.285 110.295 78.010 ;
        RECT 112.050 77.830 112.390 78.660 ;
        RECT 117.570 77.830 117.910 78.660 ;
        RECT 123.090 77.830 123.430 78.660 ;
        RECT 128.610 77.830 128.950 78.660 ;
        RECT 133.695 78.035 134.215 78.575 ;
        RECT 110.465 77.285 115.810 77.830 ;
        RECT 115.985 77.285 121.330 77.830 ;
        RECT 121.505 77.285 126.850 77.830 ;
        RECT 127.025 77.285 132.370 77.830 ;
        RECT 133.005 77.285 134.215 78.035 ;
        RECT 45.520 77.115 134.300 77.285 ;
        RECT 45.605 76.365 46.815 77.115 ;
        RECT 46.985 76.570 52.330 77.115 ;
        RECT 52.505 76.570 57.850 77.115 ;
        RECT 58.025 76.570 63.370 77.115 ;
        RECT 63.545 76.570 68.890 77.115 ;
        RECT 45.605 75.825 46.125 76.365 ;
        RECT 48.570 75.740 48.910 76.570 ;
        RECT 54.090 75.740 54.430 76.570 ;
        RECT 59.610 75.740 59.950 76.570 ;
        RECT 65.130 75.740 65.470 76.570 ;
        RECT 69.065 76.345 70.735 77.115 ;
        RECT 71.365 76.390 71.655 77.115 ;
        RECT 71.825 76.570 77.170 77.115 ;
        RECT 77.345 76.570 82.690 77.115 ;
        RECT 82.865 76.570 88.210 77.115 ;
        RECT 88.385 76.570 93.730 77.115 ;
        RECT 69.065 75.825 69.815 76.345 ;
        RECT 73.410 75.740 73.750 76.570 ;
        RECT 78.930 75.740 79.270 76.570 ;
        RECT 84.450 75.740 84.790 76.570 ;
        RECT 89.970 75.740 90.310 76.570 ;
        RECT 93.905 76.345 96.495 77.115 ;
        RECT 97.125 76.390 97.415 77.115 ;
        RECT 97.585 76.570 102.930 77.115 ;
        RECT 103.105 76.570 108.450 77.115 ;
        RECT 108.625 76.570 113.970 77.115 ;
        RECT 114.145 76.570 119.490 77.115 ;
        RECT 93.905 75.825 95.115 76.345 ;
        RECT 99.170 75.740 99.510 76.570 ;
        RECT 104.690 75.740 105.030 76.570 ;
        RECT 110.210 75.740 110.550 76.570 ;
        RECT 115.730 75.740 116.070 76.570 ;
        RECT 119.665 76.345 122.255 77.115 ;
        RECT 122.885 76.390 123.175 77.115 ;
        RECT 123.345 76.570 128.690 77.115 ;
        RECT 119.665 75.825 120.875 76.345 ;
        RECT 124.930 75.740 125.270 76.570 ;
        RECT 128.865 76.345 132.375 77.115 ;
        RECT 133.005 76.365 134.215 77.115 ;
        RECT 128.865 75.825 130.515 76.345 ;
        RECT 133.695 75.825 134.215 76.365 ;
        RECT 45.605 72.595 46.125 73.135 ;
        RECT 45.605 71.845 46.815 72.595 ;
        RECT 48.570 72.390 48.910 73.220 ;
        RECT 54.090 72.390 54.430 73.220 ;
        RECT 46.985 71.845 52.330 72.390 ;
        RECT 52.505 71.845 57.850 72.390 ;
        RECT 58.485 71.845 58.775 72.570 ;
        RECT 60.530 72.390 60.870 73.220 ;
        RECT 66.050 72.390 66.390 73.220 ;
        RECT 71.570 72.390 71.910 73.220 ;
        RECT 77.090 72.390 77.430 73.220 ;
        RECT 81.025 72.615 82.235 73.135 ;
        RECT 58.945 71.845 64.290 72.390 ;
        RECT 64.465 71.845 69.810 72.390 ;
        RECT 69.985 71.845 75.330 72.390 ;
        RECT 75.505 71.845 80.850 72.390 ;
        RECT 81.025 71.845 83.615 72.615 ;
        RECT 84.245 71.845 84.535 72.570 ;
        RECT 86.290 72.390 86.630 73.220 ;
        RECT 91.810 72.390 92.150 73.220 ;
        RECT 97.330 72.390 97.670 73.220 ;
        RECT 102.850 72.390 103.190 73.220 ;
        RECT 106.785 72.615 107.995 73.135 ;
        RECT 84.705 71.845 90.050 72.390 ;
        RECT 90.225 71.845 95.570 72.390 ;
        RECT 95.745 71.845 101.090 72.390 ;
        RECT 101.265 71.845 106.610 72.390 ;
        RECT 106.785 71.845 109.375 72.615 ;
        RECT 110.005 71.845 110.295 72.570 ;
        RECT 112.050 72.390 112.390 73.220 ;
        RECT 117.570 72.390 117.910 73.220 ;
        RECT 123.090 72.390 123.430 73.220 ;
        RECT 128.610 72.390 128.950 73.220 ;
        RECT 133.695 72.595 134.215 73.135 ;
        RECT 110.465 71.845 115.810 72.390 ;
        RECT 115.985 71.845 121.330 72.390 ;
        RECT 121.505 71.845 126.850 72.390 ;
        RECT 127.025 71.845 132.370 72.390 ;
        RECT 133.005 71.845 134.215 72.595 ;
        RECT 45.520 71.675 134.300 71.845 ;
        RECT 45.605 70.925 46.815 71.675 ;
        RECT 46.985 71.130 52.330 71.675 ;
        RECT 52.505 71.130 57.850 71.675 ;
        RECT 58.025 71.130 63.370 71.675 ;
        RECT 63.545 71.130 68.890 71.675 ;
        RECT 45.605 70.385 46.125 70.925 ;
        RECT 48.570 70.300 48.910 71.130 ;
        RECT 54.090 70.300 54.430 71.130 ;
        RECT 59.610 70.300 59.950 71.130 ;
        RECT 65.130 70.300 65.470 71.130 ;
        RECT 69.065 70.905 70.735 71.675 ;
        RECT 71.365 70.950 71.655 71.675 ;
        RECT 71.825 71.130 77.170 71.675 ;
        RECT 77.345 71.130 82.690 71.675 ;
        RECT 82.865 71.130 88.210 71.675 ;
        RECT 88.385 71.130 93.730 71.675 ;
        RECT 69.065 70.385 69.815 70.905 ;
        RECT 73.410 70.300 73.750 71.130 ;
        RECT 78.930 70.300 79.270 71.130 ;
        RECT 84.450 70.300 84.790 71.130 ;
        RECT 89.970 70.300 90.310 71.130 ;
        RECT 93.905 70.905 96.495 71.675 ;
        RECT 97.125 70.950 97.415 71.675 ;
        RECT 97.585 71.130 102.930 71.675 ;
        RECT 103.105 71.130 108.450 71.675 ;
        RECT 108.625 71.130 113.970 71.675 ;
        RECT 114.145 71.130 119.490 71.675 ;
        RECT 93.905 70.385 95.115 70.905 ;
        RECT 99.170 70.300 99.510 71.130 ;
        RECT 104.690 70.300 105.030 71.130 ;
        RECT 110.210 70.300 110.550 71.130 ;
        RECT 115.730 70.300 116.070 71.130 ;
        RECT 119.665 70.905 122.255 71.675 ;
        RECT 122.885 70.950 123.175 71.675 ;
        RECT 123.345 71.130 128.690 71.675 ;
        RECT 119.665 70.385 120.875 70.905 ;
        RECT 124.930 70.300 125.270 71.130 ;
        RECT 128.865 70.905 132.375 71.675 ;
        RECT 133.005 70.925 134.215 71.675 ;
        RECT 128.865 70.385 130.515 70.905 ;
        RECT 133.695 70.385 134.215 70.925 ;
        RECT 45.605 67.155 46.125 67.695 ;
        RECT 45.605 66.405 46.815 67.155 ;
        RECT 48.570 66.950 48.910 67.780 ;
        RECT 54.090 66.950 54.430 67.780 ;
        RECT 46.985 66.405 52.330 66.950 ;
        RECT 52.505 66.405 57.850 66.950 ;
        RECT 58.485 66.405 58.775 67.130 ;
        RECT 60.530 66.950 60.870 67.780 ;
        RECT 66.050 66.950 66.390 67.780 ;
        RECT 71.570 66.950 71.910 67.780 ;
        RECT 77.090 66.950 77.430 67.780 ;
        RECT 81.025 67.175 82.235 67.695 ;
        RECT 58.945 66.405 64.290 66.950 ;
        RECT 64.465 66.405 69.810 66.950 ;
        RECT 69.985 66.405 75.330 66.950 ;
        RECT 75.505 66.405 80.850 66.950 ;
        RECT 81.025 66.405 83.615 67.175 ;
        RECT 84.245 66.405 84.535 67.130 ;
        RECT 86.290 66.950 86.630 67.780 ;
        RECT 91.810 66.950 92.150 67.780 ;
        RECT 97.330 66.950 97.670 67.780 ;
        RECT 102.850 66.950 103.190 67.780 ;
        RECT 106.785 67.175 107.995 67.695 ;
        RECT 84.705 66.405 90.050 66.950 ;
        RECT 90.225 66.405 95.570 66.950 ;
        RECT 95.745 66.405 101.090 66.950 ;
        RECT 101.265 66.405 106.610 66.950 ;
        RECT 106.785 66.405 109.375 67.175 ;
        RECT 110.005 66.405 110.295 67.130 ;
        RECT 112.050 66.950 112.390 67.780 ;
        RECT 117.570 66.950 117.910 67.780 ;
        RECT 123.090 66.950 123.430 67.780 ;
        RECT 128.610 66.950 128.950 67.780 ;
        RECT 133.695 67.155 134.215 67.695 ;
        RECT 110.465 66.405 115.810 66.950 ;
        RECT 115.985 66.405 121.330 66.950 ;
        RECT 121.505 66.405 126.850 66.950 ;
        RECT 127.025 66.405 132.370 66.950 ;
        RECT 133.005 66.405 134.215 67.155 ;
        RECT 45.520 66.235 134.300 66.405 ;
        RECT 45.605 65.485 46.815 66.235 ;
        RECT 46.985 65.690 52.330 66.235 ;
        RECT 52.505 65.690 57.850 66.235 ;
        RECT 58.025 65.690 63.370 66.235 ;
        RECT 63.545 65.690 68.890 66.235 ;
        RECT 45.605 64.945 46.125 65.485 ;
        RECT 48.570 64.860 48.910 65.690 ;
        RECT 54.090 64.860 54.430 65.690 ;
        RECT 59.610 64.860 59.950 65.690 ;
        RECT 65.130 64.860 65.470 65.690 ;
        RECT 69.065 65.465 70.735 66.235 ;
        RECT 71.365 65.510 71.655 66.235 ;
        RECT 71.825 65.690 77.170 66.235 ;
        RECT 77.345 65.690 82.690 66.235 ;
        RECT 82.865 65.690 88.210 66.235 ;
        RECT 88.385 65.690 93.730 66.235 ;
        RECT 69.065 64.945 69.815 65.465 ;
        RECT 73.410 64.860 73.750 65.690 ;
        RECT 78.930 64.860 79.270 65.690 ;
        RECT 84.450 64.860 84.790 65.690 ;
        RECT 89.970 64.860 90.310 65.690 ;
        RECT 93.905 65.465 96.495 66.235 ;
        RECT 97.125 65.510 97.415 66.235 ;
        RECT 97.585 65.690 102.930 66.235 ;
        RECT 103.105 65.690 108.450 66.235 ;
        RECT 108.625 65.690 113.970 66.235 ;
        RECT 114.145 65.690 119.490 66.235 ;
        RECT 93.905 64.945 95.115 65.465 ;
        RECT 99.170 64.860 99.510 65.690 ;
        RECT 104.690 64.860 105.030 65.690 ;
        RECT 110.210 64.860 110.550 65.690 ;
        RECT 115.730 64.860 116.070 65.690 ;
        RECT 119.665 65.465 122.255 66.235 ;
        RECT 122.885 65.510 123.175 66.235 ;
        RECT 123.345 65.690 128.690 66.235 ;
        RECT 119.665 64.945 120.875 65.465 ;
        RECT 124.930 64.860 125.270 65.690 ;
        RECT 128.865 65.465 132.375 66.235 ;
        RECT 133.005 65.485 134.215 66.235 ;
        RECT 128.865 64.945 130.515 65.465 ;
        RECT 133.695 64.945 134.215 65.485 ;
        RECT 45.605 61.715 46.125 62.255 ;
        RECT 45.605 60.965 46.815 61.715 ;
        RECT 48.570 61.510 48.910 62.340 ;
        RECT 54.090 61.510 54.430 62.340 ;
        RECT 46.985 60.965 52.330 61.510 ;
        RECT 52.505 60.965 57.850 61.510 ;
        RECT 58.485 60.965 58.775 61.690 ;
        RECT 60.530 61.510 60.870 62.340 ;
        RECT 66.050 61.510 66.390 62.340 ;
        RECT 69.985 61.715 70.505 62.255 ;
        RECT 58.945 60.965 64.290 61.510 ;
        RECT 64.465 60.965 69.810 61.510 ;
        RECT 69.985 60.965 71.195 61.715 ;
        RECT 71.365 60.965 71.655 61.690 ;
        RECT 73.410 61.510 73.750 62.340 ;
        RECT 78.930 61.510 79.270 62.340 ;
        RECT 82.865 61.715 83.385 62.255 ;
        RECT 71.825 60.965 77.170 61.510 ;
        RECT 77.345 60.965 82.690 61.510 ;
        RECT 82.865 60.965 84.075 61.715 ;
        RECT 84.245 60.965 84.535 61.690 ;
        RECT 86.290 61.510 86.630 62.340 ;
        RECT 91.810 61.510 92.150 62.340 ;
        RECT 95.745 61.715 96.265 62.255 ;
        RECT 84.705 60.965 90.050 61.510 ;
        RECT 90.225 60.965 95.570 61.510 ;
        RECT 95.745 60.965 96.955 61.715 ;
        RECT 97.125 60.965 97.415 61.690 ;
        RECT 99.170 61.510 99.510 62.340 ;
        RECT 104.690 61.510 105.030 62.340 ;
        RECT 108.625 61.715 109.145 62.255 ;
        RECT 97.585 60.965 102.930 61.510 ;
        RECT 103.105 60.965 108.450 61.510 ;
        RECT 108.625 60.965 109.835 61.715 ;
        RECT 110.005 60.965 110.295 61.690 ;
        RECT 112.050 61.510 112.390 62.340 ;
        RECT 117.570 61.510 117.910 62.340 ;
        RECT 121.505 61.715 122.025 62.255 ;
        RECT 110.465 60.965 115.810 61.510 ;
        RECT 115.985 60.965 121.330 61.510 ;
        RECT 121.505 60.965 122.715 61.715 ;
        RECT 122.885 60.965 123.175 61.690 ;
        RECT 124.930 61.510 125.270 62.340 ;
        RECT 128.865 61.735 130.515 62.255 ;
        RECT 123.345 60.965 128.690 61.510 ;
        RECT 128.865 60.965 132.375 61.735 ;
        RECT 133.695 61.715 134.215 62.255 ;
        RECT 133.005 60.965 134.215 61.715 ;
        RECT 45.520 60.795 134.300 60.965 ;
      LAYER mcon ;
        RECT 45.665 136.955 45.835 137.125 ;
        RECT 46.125 136.955 46.295 137.125 ;
        RECT 46.585 136.955 46.755 137.125 ;
        RECT 47.045 136.955 47.215 137.125 ;
        RECT 47.505 136.955 47.675 137.125 ;
        RECT 47.965 136.955 48.135 137.125 ;
        RECT 48.425 136.955 48.595 137.125 ;
        RECT 48.885 136.955 49.055 137.125 ;
        RECT 49.345 136.955 49.515 137.125 ;
        RECT 49.805 136.955 49.975 137.125 ;
        RECT 50.265 136.955 50.435 137.125 ;
        RECT 50.725 136.955 50.895 137.125 ;
        RECT 51.185 136.955 51.355 137.125 ;
        RECT 51.645 136.955 51.815 137.125 ;
        RECT 52.105 136.955 52.275 137.125 ;
        RECT 52.565 136.955 52.735 137.125 ;
        RECT 53.025 136.955 53.195 137.125 ;
        RECT 53.485 136.955 53.655 137.125 ;
        RECT 53.945 136.955 54.115 137.125 ;
        RECT 54.405 136.955 54.575 137.125 ;
        RECT 54.865 136.955 55.035 137.125 ;
        RECT 55.325 136.955 55.495 137.125 ;
        RECT 55.785 136.955 55.955 137.125 ;
        RECT 56.245 136.955 56.415 137.125 ;
        RECT 56.705 136.955 56.875 137.125 ;
        RECT 57.165 136.955 57.335 137.125 ;
        RECT 57.625 136.955 57.795 137.125 ;
        RECT 58.085 136.955 58.255 137.125 ;
        RECT 58.545 136.955 58.715 137.125 ;
        RECT 59.005 136.955 59.175 137.125 ;
        RECT 59.465 136.955 59.635 137.125 ;
        RECT 59.925 136.955 60.095 137.125 ;
        RECT 60.385 136.955 60.555 137.125 ;
        RECT 60.845 136.955 61.015 137.125 ;
        RECT 61.305 136.955 61.475 137.125 ;
        RECT 61.765 136.955 61.935 137.125 ;
        RECT 62.225 136.955 62.395 137.125 ;
        RECT 62.685 136.955 62.855 137.125 ;
        RECT 63.145 136.955 63.315 137.125 ;
        RECT 63.605 136.955 63.775 137.125 ;
        RECT 64.065 136.955 64.235 137.125 ;
        RECT 64.525 136.955 64.695 137.125 ;
        RECT 64.985 136.955 65.155 137.125 ;
        RECT 65.445 136.955 65.615 137.125 ;
        RECT 65.905 136.955 66.075 137.125 ;
        RECT 66.365 136.955 66.535 137.125 ;
        RECT 66.825 136.955 66.995 137.125 ;
        RECT 67.285 136.955 67.455 137.125 ;
        RECT 67.745 136.955 67.915 137.125 ;
        RECT 68.205 136.955 68.375 137.125 ;
        RECT 68.665 136.955 68.835 137.125 ;
        RECT 69.125 136.955 69.295 137.125 ;
        RECT 69.585 136.955 69.755 137.125 ;
        RECT 70.045 136.955 70.215 137.125 ;
        RECT 70.505 136.955 70.675 137.125 ;
        RECT 70.965 136.955 71.135 137.125 ;
        RECT 71.425 136.955 71.595 137.125 ;
        RECT 71.885 136.955 72.055 137.125 ;
        RECT 72.345 136.955 72.515 137.125 ;
        RECT 72.805 136.955 72.975 137.125 ;
        RECT 73.265 136.955 73.435 137.125 ;
        RECT 73.725 136.955 73.895 137.125 ;
        RECT 74.185 136.955 74.355 137.125 ;
        RECT 74.645 136.955 74.815 137.125 ;
        RECT 75.105 136.955 75.275 137.125 ;
        RECT 75.565 136.955 75.735 137.125 ;
        RECT 76.025 136.955 76.195 137.125 ;
        RECT 76.485 136.955 76.655 137.125 ;
        RECT 76.945 136.955 77.115 137.125 ;
        RECT 77.405 136.955 77.575 137.125 ;
        RECT 77.865 136.955 78.035 137.125 ;
        RECT 78.325 136.955 78.495 137.125 ;
        RECT 78.785 136.955 78.955 137.125 ;
        RECT 79.245 136.955 79.415 137.125 ;
        RECT 79.705 136.955 79.875 137.125 ;
        RECT 80.165 136.955 80.335 137.125 ;
        RECT 80.625 136.955 80.795 137.125 ;
        RECT 81.085 136.955 81.255 137.125 ;
        RECT 81.545 136.955 81.715 137.125 ;
        RECT 82.005 136.955 82.175 137.125 ;
        RECT 82.465 136.955 82.635 137.125 ;
        RECT 82.925 136.955 83.095 137.125 ;
        RECT 83.385 136.955 83.555 137.125 ;
        RECT 83.845 136.955 84.015 137.125 ;
        RECT 84.305 136.955 84.475 137.125 ;
        RECT 84.765 136.955 84.935 137.125 ;
        RECT 85.225 136.955 85.395 137.125 ;
        RECT 85.685 136.955 85.855 137.125 ;
        RECT 86.145 136.955 86.315 137.125 ;
        RECT 86.605 136.955 86.775 137.125 ;
        RECT 87.065 136.955 87.235 137.125 ;
        RECT 87.525 136.955 87.695 137.125 ;
        RECT 87.985 136.955 88.155 137.125 ;
        RECT 88.445 136.955 88.615 137.125 ;
        RECT 88.905 136.955 89.075 137.125 ;
        RECT 89.365 136.955 89.535 137.125 ;
        RECT 89.825 136.955 89.995 137.125 ;
        RECT 90.285 136.955 90.455 137.125 ;
        RECT 90.745 136.955 90.915 137.125 ;
        RECT 91.205 136.955 91.375 137.125 ;
        RECT 91.665 136.955 91.835 137.125 ;
        RECT 92.125 136.955 92.295 137.125 ;
        RECT 92.585 136.955 92.755 137.125 ;
        RECT 93.045 136.955 93.215 137.125 ;
        RECT 93.505 136.955 93.675 137.125 ;
        RECT 93.965 136.955 94.135 137.125 ;
        RECT 94.425 136.955 94.595 137.125 ;
        RECT 94.885 136.955 95.055 137.125 ;
        RECT 95.345 136.955 95.515 137.125 ;
        RECT 95.805 136.955 95.975 137.125 ;
        RECT 96.265 136.955 96.435 137.125 ;
        RECT 96.725 136.955 96.895 137.125 ;
        RECT 97.185 136.955 97.355 137.125 ;
        RECT 97.645 136.955 97.815 137.125 ;
        RECT 98.105 136.955 98.275 137.125 ;
        RECT 98.565 136.955 98.735 137.125 ;
        RECT 99.025 136.955 99.195 137.125 ;
        RECT 99.485 136.955 99.655 137.125 ;
        RECT 99.945 136.955 100.115 137.125 ;
        RECT 100.405 136.955 100.575 137.125 ;
        RECT 100.865 136.955 101.035 137.125 ;
        RECT 101.325 136.955 101.495 137.125 ;
        RECT 101.785 136.955 101.955 137.125 ;
        RECT 102.245 136.955 102.415 137.125 ;
        RECT 102.705 136.955 102.875 137.125 ;
        RECT 103.165 136.955 103.335 137.125 ;
        RECT 103.625 136.955 103.795 137.125 ;
        RECT 104.085 136.955 104.255 137.125 ;
        RECT 104.545 136.955 104.715 137.125 ;
        RECT 105.005 136.955 105.175 137.125 ;
        RECT 105.465 136.955 105.635 137.125 ;
        RECT 105.925 136.955 106.095 137.125 ;
        RECT 106.385 136.955 106.555 137.125 ;
        RECT 106.845 136.955 107.015 137.125 ;
        RECT 107.305 136.955 107.475 137.125 ;
        RECT 107.765 136.955 107.935 137.125 ;
        RECT 108.225 136.955 108.395 137.125 ;
        RECT 108.685 136.955 108.855 137.125 ;
        RECT 109.145 136.955 109.315 137.125 ;
        RECT 109.605 136.955 109.775 137.125 ;
        RECT 110.065 136.955 110.235 137.125 ;
        RECT 110.525 136.955 110.695 137.125 ;
        RECT 110.985 136.955 111.155 137.125 ;
        RECT 111.445 136.955 111.615 137.125 ;
        RECT 111.905 136.955 112.075 137.125 ;
        RECT 112.365 136.955 112.535 137.125 ;
        RECT 112.825 136.955 112.995 137.125 ;
        RECT 113.285 136.955 113.455 137.125 ;
        RECT 113.745 136.955 113.915 137.125 ;
        RECT 114.205 136.955 114.375 137.125 ;
        RECT 114.665 136.955 114.835 137.125 ;
        RECT 115.125 136.955 115.295 137.125 ;
        RECT 115.585 136.955 115.755 137.125 ;
        RECT 116.045 136.955 116.215 137.125 ;
        RECT 116.505 136.955 116.675 137.125 ;
        RECT 116.965 136.955 117.135 137.125 ;
        RECT 117.425 136.955 117.595 137.125 ;
        RECT 117.885 136.955 118.055 137.125 ;
        RECT 118.345 136.955 118.515 137.125 ;
        RECT 118.805 136.955 118.975 137.125 ;
        RECT 119.265 136.955 119.435 137.125 ;
        RECT 119.725 136.955 119.895 137.125 ;
        RECT 120.185 136.955 120.355 137.125 ;
        RECT 120.645 136.955 120.815 137.125 ;
        RECT 121.105 136.955 121.275 137.125 ;
        RECT 121.565 136.955 121.735 137.125 ;
        RECT 122.025 136.955 122.195 137.125 ;
        RECT 122.485 136.955 122.655 137.125 ;
        RECT 122.945 136.955 123.115 137.125 ;
        RECT 123.405 136.955 123.575 137.125 ;
        RECT 123.865 136.955 124.035 137.125 ;
        RECT 124.325 136.955 124.495 137.125 ;
        RECT 124.785 136.955 124.955 137.125 ;
        RECT 125.245 136.955 125.415 137.125 ;
        RECT 125.705 136.955 125.875 137.125 ;
        RECT 126.165 136.955 126.335 137.125 ;
        RECT 126.625 136.955 126.795 137.125 ;
        RECT 127.085 136.955 127.255 137.125 ;
        RECT 127.545 136.955 127.715 137.125 ;
        RECT 128.005 136.955 128.175 137.125 ;
        RECT 128.465 136.955 128.635 137.125 ;
        RECT 128.925 136.955 129.095 137.125 ;
        RECT 129.385 136.955 129.555 137.125 ;
        RECT 129.845 136.955 130.015 137.125 ;
        RECT 130.305 136.955 130.475 137.125 ;
        RECT 130.765 136.955 130.935 137.125 ;
        RECT 131.225 136.955 131.395 137.125 ;
        RECT 131.685 136.955 131.855 137.125 ;
        RECT 132.145 136.955 132.315 137.125 ;
        RECT 132.605 136.955 132.775 137.125 ;
        RECT 133.065 136.955 133.235 137.125 ;
        RECT 133.525 136.955 133.695 137.125 ;
        RECT 133.985 136.955 134.155 137.125 ;
        RECT 45.665 131.515 45.835 131.685 ;
        RECT 46.125 131.515 46.295 131.685 ;
        RECT 46.585 131.515 46.755 131.685 ;
        RECT 47.045 131.515 47.215 131.685 ;
        RECT 47.505 131.515 47.675 131.685 ;
        RECT 47.965 131.515 48.135 131.685 ;
        RECT 48.425 131.515 48.595 131.685 ;
        RECT 48.885 131.515 49.055 131.685 ;
        RECT 49.345 131.515 49.515 131.685 ;
        RECT 49.805 131.515 49.975 131.685 ;
        RECT 50.265 131.515 50.435 131.685 ;
        RECT 50.725 131.515 50.895 131.685 ;
        RECT 51.185 131.515 51.355 131.685 ;
        RECT 51.645 131.515 51.815 131.685 ;
        RECT 52.105 131.515 52.275 131.685 ;
        RECT 52.565 131.515 52.735 131.685 ;
        RECT 53.025 131.515 53.195 131.685 ;
        RECT 53.485 131.515 53.655 131.685 ;
        RECT 53.945 131.515 54.115 131.685 ;
        RECT 54.405 131.515 54.575 131.685 ;
        RECT 54.865 131.515 55.035 131.685 ;
        RECT 55.325 131.515 55.495 131.685 ;
        RECT 55.785 131.515 55.955 131.685 ;
        RECT 56.245 131.515 56.415 131.685 ;
        RECT 56.705 131.515 56.875 131.685 ;
        RECT 57.165 131.515 57.335 131.685 ;
        RECT 57.625 131.515 57.795 131.685 ;
        RECT 58.085 131.515 58.255 131.685 ;
        RECT 58.545 131.515 58.715 131.685 ;
        RECT 59.005 131.515 59.175 131.685 ;
        RECT 59.465 131.515 59.635 131.685 ;
        RECT 59.925 131.515 60.095 131.685 ;
        RECT 60.385 131.515 60.555 131.685 ;
        RECT 60.845 131.515 61.015 131.685 ;
        RECT 61.305 131.515 61.475 131.685 ;
        RECT 61.765 131.515 61.935 131.685 ;
        RECT 62.225 131.515 62.395 131.685 ;
        RECT 62.685 131.515 62.855 131.685 ;
        RECT 63.145 131.515 63.315 131.685 ;
        RECT 63.605 131.515 63.775 131.685 ;
        RECT 64.065 131.515 64.235 131.685 ;
        RECT 64.525 131.515 64.695 131.685 ;
        RECT 64.985 131.515 65.155 131.685 ;
        RECT 65.445 131.515 65.615 131.685 ;
        RECT 65.905 131.515 66.075 131.685 ;
        RECT 66.365 131.515 66.535 131.685 ;
        RECT 66.825 131.515 66.995 131.685 ;
        RECT 67.285 131.515 67.455 131.685 ;
        RECT 67.745 131.515 67.915 131.685 ;
        RECT 68.205 131.515 68.375 131.685 ;
        RECT 68.665 131.515 68.835 131.685 ;
        RECT 69.125 131.515 69.295 131.685 ;
        RECT 69.585 131.515 69.755 131.685 ;
        RECT 70.045 131.515 70.215 131.685 ;
        RECT 70.505 131.515 70.675 131.685 ;
        RECT 70.965 131.515 71.135 131.685 ;
        RECT 71.425 131.515 71.595 131.685 ;
        RECT 71.885 131.515 72.055 131.685 ;
        RECT 72.345 131.515 72.515 131.685 ;
        RECT 72.805 131.515 72.975 131.685 ;
        RECT 73.265 131.515 73.435 131.685 ;
        RECT 73.725 131.515 73.895 131.685 ;
        RECT 74.185 131.515 74.355 131.685 ;
        RECT 74.645 131.515 74.815 131.685 ;
        RECT 75.105 131.515 75.275 131.685 ;
        RECT 75.565 131.515 75.735 131.685 ;
        RECT 76.025 131.515 76.195 131.685 ;
        RECT 76.485 131.515 76.655 131.685 ;
        RECT 76.945 131.515 77.115 131.685 ;
        RECT 77.405 131.515 77.575 131.685 ;
        RECT 77.865 131.515 78.035 131.685 ;
        RECT 78.325 131.515 78.495 131.685 ;
        RECT 78.785 131.515 78.955 131.685 ;
        RECT 79.245 131.515 79.415 131.685 ;
        RECT 79.705 131.515 79.875 131.685 ;
        RECT 80.165 131.515 80.335 131.685 ;
        RECT 80.625 131.515 80.795 131.685 ;
        RECT 81.085 131.515 81.255 131.685 ;
        RECT 81.545 131.515 81.715 131.685 ;
        RECT 82.005 131.515 82.175 131.685 ;
        RECT 82.465 131.515 82.635 131.685 ;
        RECT 82.925 131.515 83.095 131.685 ;
        RECT 83.385 131.515 83.555 131.685 ;
        RECT 83.845 131.515 84.015 131.685 ;
        RECT 84.305 131.515 84.475 131.685 ;
        RECT 84.765 131.515 84.935 131.685 ;
        RECT 85.225 131.515 85.395 131.685 ;
        RECT 85.685 131.515 85.855 131.685 ;
        RECT 86.145 131.515 86.315 131.685 ;
        RECT 86.605 131.515 86.775 131.685 ;
        RECT 87.065 131.515 87.235 131.685 ;
        RECT 87.525 131.515 87.695 131.685 ;
        RECT 87.985 131.515 88.155 131.685 ;
        RECT 88.445 131.515 88.615 131.685 ;
        RECT 88.905 131.515 89.075 131.685 ;
        RECT 89.365 131.515 89.535 131.685 ;
        RECT 89.825 131.515 89.995 131.685 ;
        RECT 90.285 131.515 90.455 131.685 ;
        RECT 90.745 131.515 90.915 131.685 ;
        RECT 91.205 131.515 91.375 131.685 ;
        RECT 91.665 131.515 91.835 131.685 ;
        RECT 92.125 131.515 92.295 131.685 ;
        RECT 92.585 131.515 92.755 131.685 ;
        RECT 93.045 131.515 93.215 131.685 ;
        RECT 93.505 131.515 93.675 131.685 ;
        RECT 93.965 131.515 94.135 131.685 ;
        RECT 94.425 131.515 94.595 131.685 ;
        RECT 94.885 131.515 95.055 131.685 ;
        RECT 95.345 131.515 95.515 131.685 ;
        RECT 95.805 131.515 95.975 131.685 ;
        RECT 96.265 131.515 96.435 131.685 ;
        RECT 96.725 131.515 96.895 131.685 ;
        RECT 97.185 131.515 97.355 131.685 ;
        RECT 97.645 131.515 97.815 131.685 ;
        RECT 98.105 131.515 98.275 131.685 ;
        RECT 98.565 131.515 98.735 131.685 ;
        RECT 99.025 131.515 99.195 131.685 ;
        RECT 99.485 131.515 99.655 131.685 ;
        RECT 99.945 131.515 100.115 131.685 ;
        RECT 100.405 131.515 100.575 131.685 ;
        RECT 100.865 131.515 101.035 131.685 ;
        RECT 101.325 131.515 101.495 131.685 ;
        RECT 101.785 131.515 101.955 131.685 ;
        RECT 102.245 131.515 102.415 131.685 ;
        RECT 102.705 131.515 102.875 131.685 ;
        RECT 103.165 131.515 103.335 131.685 ;
        RECT 103.625 131.515 103.795 131.685 ;
        RECT 104.085 131.515 104.255 131.685 ;
        RECT 104.545 131.515 104.715 131.685 ;
        RECT 105.005 131.515 105.175 131.685 ;
        RECT 105.465 131.515 105.635 131.685 ;
        RECT 105.925 131.515 106.095 131.685 ;
        RECT 106.385 131.515 106.555 131.685 ;
        RECT 106.845 131.515 107.015 131.685 ;
        RECT 107.305 131.515 107.475 131.685 ;
        RECT 107.765 131.515 107.935 131.685 ;
        RECT 108.225 131.515 108.395 131.685 ;
        RECT 108.685 131.515 108.855 131.685 ;
        RECT 109.145 131.515 109.315 131.685 ;
        RECT 109.605 131.515 109.775 131.685 ;
        RECT 110.065 131.515 110.235 131.685 ;
        RECT 110.525 131.515 110.695 131.685 ;
        RECT 110.985 131.515 111.155 131.685 ;
        RECT 111.445 131.515 111.615 131.685 ;
        RECT 111.905 131.515 112.075 131.685 ;
        RECT 112.365 131.515 112.535 131.685 ;
        RECT 112.825 131.515 112.995 131.685 ;
        RECT 113.285 131.515 113.455 131.685 ;
        RECT 113.745 131.515 113.915 131.685 ;
        RECT 114.205 131.515 114.375 131.685 ;
        RECT 114.665 131.515 114.835 131.685 ;
        RECT 115.125 131.515 115.295 131.685 ;
        RECT 115.585 131.515 115.755 131.685 ;
        RECT 116.045 131.515 116.215 131.685 ;
        RECT 116.505 131.515 116.675 131.685 ;
        RECT 116.965 131.515 117.135 131.685 ;
        RECT 117.425 131.515 117.595 131.685 ;
        RECT 117.885 131.515 118.055 131.685 ;
        RECT 118.345 131.515 118.515 131.685 ;
        RECT 118.805 131.515 118.975 131.685 ;
        RECT 119.265 131.515 119.435 131.685 ;
        RECT 119.725 131.515 119.895 131.685 ;
        RECT 120.185 131.515 120.355 131.685 ;
        RECT 120.645 131.515 120.815 131.685 ;
        RECT 121.105 131.515 121.275 131.685 ;
        RECT 121.565 131.515 121.735 131.685 ;
        RECT 122.025 131.515 122.195 131.685 ;
        RECT 122.485 131.515 122.655 131.685 ;
        RECT 122.945 131.515 123.115 131.685 ;
        RECT 123.405 131.515 123.575 131.685 ;
        RECT 123.865 131.515 124.035 131.685 ;
        RECT 124.325 131.515 124.495 131.685 ;
        RECT 124.785 131.515 124.955 131.685 ;
        RECT 125.245 131.515 125.415 131.685 ;
        RECT 125.705 131.515 125.875 131.685 ;
        RECT 126.165 131.515 126.335 131.685 ;
        RECT 126.625 131.515 126.795 131.685 ;
        RECT 127.085 131.515 127.255 131.685 ;
        RECT 127.545 131.515 127.715 131.685 ;
        RECT 128.005 131.515 128.175 131.685 ;
        RECT 128.465 131.515 128.635 131.685 ;
        RECT 128.925 131.515 129.095 131.685 ;
        RECT 129.385 131.515 129.555 131.685 ;
        RECT 129.845 131.515 130.015 131.685 ;
        RECT 130.305 131.515 130.475 131.685 ;
        RECT 130.765 131.515 130.935 131.685 ;
        RECT 131.225 131.515 131.395 131.685 ;
        RECT 131.685 131.515 131.855 131.685 ;
        RECT 132.145 131.515 132.315 131.685 ;
        RECT 132.605 131.515 132.775 131.685 ;
        RECT 133.065 131.515 133.235 131.685 ;
        RECT 133.525 131.515 133.695 131.685 ;
        RECT 133.985 131.515 134.155 131.685 ;
        RECT 45.665 126.075 45.835 126.245 ;
        RECT 46.125 126.075 46.295 126.245 ;
        RECT 46.585 126.075 46.755 126.245 ;
        RECT 47.045 126.075 47.215 126.245 ;
        RECT 47.505 126.075 47.675 126.245 ;
        RECT 47.965 126.075 48.135 126.245 ;
        RECT 48.425 126.075 48.595 126.245 ;
        RECT 48.885 126.075 49.055 126.245 ;
        RECT 49.345 126.075 49.515 126.245 ;
        RECT 49.805 126.075 49.975 126.245 ;
        RECT 50.265 126.075 50.435 126.245 ;
        RECT 50.725 126.075 50.895 126.245 ;
        RECT 51.185 126.075 51.355 126.245 ;
        RECT 51.645 126.075 51.815 126.245 ;
        RECT 52.105 126.075 52.275 126.245 ;
        RECT 52.565 126.075 52.735 126.245 ;
        RECT 53.025 126.075 53.195 126.245 ;
        RECT 53.485 126.075 53.655 126.245 ;
        RECT 53.945 126.075 54.115 126.245 ;
        RECT 54.405 126.075 54.575 126.245 ;
        RECT 54.865 126.075 55.035 126.245 ;
        RECT 55.325 126.075 55.495 126.245 ;
        RECT 55.785 126.075 55.955 126.245 ;
        RECT 56.245 126.075 56.415 126.245 ;
        RECT 56.705 126.075 56.875 126.245 ;
        RECT 57.165 126.075 57.335 126.245 ;
        RECT 57.625 126.075 57.795 126.245 ;
        RECT 58.085 126.075 58.255 126.245 ;
        RECT 58.545 126.075 58.715 126.245 ;
        RECT 59.005 126.075 59.175 126.245 ;
        RECT 59.465 126.075 59.635 126.245 ;
        RECT 59.925 126.075 60.095 126.245 ;
        RECT 60.385 126.075 60.555 126.245 ;
        RECT 60.845 126.075 61.015 126.245 ;
        RECT 61.305 126.075 61.475 126.245 ;
        RECT 61.765 126.075 61.935 126.245 ;
        RECT 62.225 126.075 62.395 126.245 ;
        RECT 62.685 126.075 62.855 126.245 ;
        RECT 63.145 126.075 63.315 126.245 ;
        RECT 63.605 126.075 63.775 126.245 ;
        RECT 64.065 126.075 64.235 126.245 ;
        RECT 64.525 126.075 64.695 126.245 ;
        RECT 64.985 126.075 65.155 126.245 ;
        RECT 65.445 126.075 65.615 126.245 ;
        RECT 65.905 126.075 66.075 126.245 ;
        RECT 66.365 126.075 66.535 126.245 ;
        RECT 66.825 126.075 66.995 126.245 ;
        RECT 67.285 126.075 67.455 126.245 ;
        RECT 67.745 126.075 67.915 126.245 ;
        RECT 68.205 126.075 68.375 126.245 ;
        RECT 68.665 126.075 68.835 126.245 ;
        RECT 69.125 126.075 69.295 126.245 ;
        RECT 69.585 126.075 69.755 126.245 ;
        RECT 70.045 126.075 70.215 126.245 ;
        RECT 70.505 126.075 70.675 126.245 ;
        RECT 70.965 126.075 71.135 126.245 ;
        RECT 71.425 126.075 71.595 126.245 ;
        RECT 71.885 126.075 72.055 126.245 ;
        RECT 72.345 126.075 72.515 126.245 ;
        RECT 72.805 126.075 72.975 126.245 ;
        RECT 73.265 126.075 73.435 126.245 ;
        RECT 73.725 126.075 73.895 126.245 ;
        RECT 74.185 126.075 74.355 126.245 ;
        RECT 74.645 126.075 74.815 126.245 ;
        RECT 75.105 126.075 75.275 126.245 ;
        RECT 75.565 126.075 75.735 126.245 ;
        RECT 76.025 126.075 76.195 126.245 ;
        RECT 76.485 126.075 76.655 126.245 ;
        RECT 76.945 126.075 77.115 126.245 ;
        RECT 77.405 126.075 77.575 126.245 ;
        RECT 77.865 126.075 78.035 126.245 ;
        RECT 78.325 126.075 78.495 126.245 ;
        RECT 78.785 126.075 78.955 126.245 ;
        RECT 79.245 126.075 79.415 126.245 ;
        RECT 79.705 126.075 79.875 126.245 ;
        RECT 80.165 126.075 80.335 126.245 ;
        RECT 80.625 126.075 80.795 126.245 ;
        RECT 81.085 126.075 81.255 126.245 ;
        RECT 81.545 126.075 81.715 126.245 ;
        RECT 82.005 126.075 82.175 126.245 ;
        RECT 82.465 126.075 82.635 126.245 ;
        RECT 82.925 126.075 83.095 126.245 ;
        RECT 83.385 126.075 83.555 126.245 ;
        RECT 83.845 126.075 84.015 126.245 ;
        RECT 84.305 126.075 84.475 126.245 ;
        RECT 84.765 126.075 84.935 126.245 ;
        RECT 85.225 126.075 85.395 126.245 ;
        RECT 85.685 126.075 85.855 126.245 ;
        RECT 86.145 126.075 86.315 126.245 ;
        RECT 86.605 126.075 86.775 126.245 ;
        RECT 87.065 126.075 87.235 126.245 ;
        RECT 87.525 126.075 87.695 126.245 ;
        RECT 87.985 126.075 88.155 126.245 ;
        RECT 88.445 126.075 88.615 126.245 ;
        RECT 88.905 126.075 89.075 126.245 ;
        RECT 89.365 126.075 89.535 126.245 ;
        RECT 89.825 126.075 89.995 126.245 ;
        RECT 90.285 126.075 90.455 126.245 ;
        RECT 90.745 126.075 90.915 126.245 ;
        RECT 91.205 126.075 91.375 126.245 ;
        RECT 91.665 126.075 91.835 126.245 ;
        RECT 92.125 126.075 92.295 126.245 ;
        RECT 92.585 126.075 92.755 126.245 ;
        RECT 93.045 126.075 93.215 126.245 ;
        RECT 93.505 126.075 93.675 126.245 ;
        RECT 93.965 126.075 94.135 126.245 ;
        RECT 94.425 126.075 94.595 126.245 ;
        RECT 94.885 126.075 95.055 126.245 ;
        RECT 95.345 126.075 95.515 126.245 ;
        RECT 95.805 126.075 95.975 126.245 ;
        RECT 96.265 126.075 96.435 126.245 ;
        RECT 96.725 126.075 96.895 126.245 ;
        RECT 97.185 126.075 97.355 126.245 ;
        RECT 97.645 126.075 97.815 126.245 ;
        RECT 98.105 126.075 98.275 126.245 ;
        RECT 98.565 126.075 98.735 126.245 ;
        RECT 99.025 126.075 99.195 126.245 ;
        RECT 99.485 126.075 99.655 126.245 ;
        RECT 99.945 126.075 100.115 126.245 ;
        RECT 100.405 126.075 100.575 126.245 ;
        RECT 100.865 126.075 101.035 126.245 ;
        RECT 101.325 126.075 101.495 126.245 ;
        RECT 101.785 126.075 101.955 126.245 ;
        RECT 102.245 126.075 102.415 126.245 ;
        RECT 102.705 126.075 102.875 126.245 ;
        RECT 103.165 126.075 103.335 126.245 ;
        RECT 103.625 126.075 103.795 126.245 ;
        RECT 104.085 126.075 104.255 126.245 ;
        RECT 104.545 126.075 104.715 126.245 ;
        RECT 105.005 126.075 105.175 126.245 ;
        RECT 105.465 126.075 105.635 126.245 ;
        RECT 105.925 126.075 106.095 126.245 ;
        RECT 106.385 126.075 106.555 126.245 ;
        RECT 106.845 126.075 107.015 126.245 ;
        RECT 107.305 126.075 107.475 126.245 ;
        RECT 107.765 126.075 107.935 126.245 ;
        RECT 108.225 126.075 108.395 126.245 ;
        RECT 108.685 126.075 108.855 126.245 ;
        RECT 109.145 126.075 109.315 126.245 ;
        RECT 109.605 126.075 109.775 126.245 ;
        RECT 110.065 126.075 110.235 126.245 ;
        RECT 110.525 126.075 110.695 126.245 ;
        RECT 110.985 126.075 111.155 126.245 ;
        RECT 111.445 126.075 111.615 126.245 ;
        RECT 111.905 126.075 112.075 126.245 ;
        RECT 112.365 126.075 112.535 126.245 ;
        RECT 112.825 126.075 112.995 126.245 ;
        RECT 113.285 126.075 113.455 126.245 ;
        RECT 113.745 126.075 113.915 126.245 ;
        RECT 114.205 126.075 114.375 126.245 ;
        RECT 114.665 126.075 114.835 126.245 ;
        RECT 115.125 126.075 115.295 126.245 ;
        RECT 115.585 126.075 115.755 126.245 ;
        RECT 116.045 126.075 116.215 126.245 ;
        RECT 116.505 126.075 116.675 126.245 ;
        RECT 116.965 126.075 117.135 126.245 ;
        RECT 117.425 126.075 117.595 126.245 ;
        RECT 117.885 126.075 118.055 126.245 ;
        RECT 118.345 126.075 118.515 126.245 ;
        RECT 118.805 126.075 118.975 126.245 ;
        RECT 119.265 126.075 119.435 126.245 ;
        RECT 119.725 126.075 119.895 126.245 ;
        RECT 120.185 126.075 120.355 126.245 ;
        RECT 120.645 126.075 120.815 126.245 ;
        RECT 121.105 126.075 121.275 126.245 ;
        RECT 121.565 126.075 121.735 126.245 ;
        RECT 122.025 126.075 122.195 126.245 ;
        RECT 122.485 126.075 122.655 126.245 ;
        RECT 122.945 126.075 123.115 126.245 ;
        RECT 123.405 126.075 123.575 126.245 ;
        RECT 123.865 126.075 124.035 126.245 ;
        RECT 124.325 126.075 124.495 126.245 ;
        RECT 124.785 126.075 124.955 126.245 ;
        RECT 125.245 126.075 125.415 126.245 ;
        RECT 125.705 126.075 125.875 126.245 ;
        RECT 126.165 126.075 126.335 126.245 ;
        RECT 126.625 126.075 126.795 126.245 ;
        RECT 127.085 126.075 127.255 126.245 ;
        RECT 127.545 126.075 127.715 126.245 ;
        RECT 128.005 126.075 128.175 126.245 ;
        RECT 128.465 126.075 128.635 126.245 ;
        RECT 128.925 126.075 129.095 126.245 ;
        RECT 129.385 126.075 129.555 126.245 ;
        RECT 129.845 126.075 130.015 126.245 ;
        RECT 130.305 126.075 130.475 126.245 ;
        RECT 130.765 126.075 130.935 126.245 ;
        RECT 131.225 126.075 131.395 126.245 ;
        RECT 131.685 126.075 131.855 126.245 ;
        RECT 132.145 126.075 132.315 126.245 ;
        RECT 132.605 126.075 132.775 126.245 ;
        RECT 133.065 126.075 133.235 126.245 ;
        RECT 133.525 126.075 133.695 126.245 ;
        RECT 133.985 126.075 134.155 126.245 ;
        RECT 45.665 120.635 45.835 120.805 ;
        RECT 46.125 120.635 46.295 120.805 ;
        RECT 46.585 120.635 46.755 120.805 ;
        RECT 47.045 120.635 47.215 120.805 ;
        RECT 47.505 120.635 47.675 120.805 ;
        RECT 47.965 120.635 48.135 120.805 ;
        RECT 48.425 120.635 48.595 120.805 ;
        RECT 48.885 120.635 49.055 120.805 ;
        RECT 49.345 120.635 49.515 120.805 ;
        RECT 49.805 120.635 49.975 120.805 ;
        RECT 50.265 120.635 50.435 120.805 ;
        RECT 50.725 120.635 50.895 120.805 ;
        RECT 51.185 120.635 51.355 120.805 ;
        RECT 51.645 120.635 51.815 120.805 ;
        RECT 52.105 120.635 52.275 120.805 ;
        RECT 52.565 120.635 52.735 120.805 ;
        RECT 53.025 120.635 53.195 120.805 ;
        RECT 53.485 120.635 53.655 120.805 ;
        RECT 53.945 120.635 54.115 120.805 ;
        RECT 54.405 120.635 54.575 120.805 ;
        RECT 54.865 120.635 55.035 120.805 ;
        RECT 55.325 120.635 55.495 120.805 ;
        RECT 55.785 120.635 55.955 120.805 ;
        RECT 56.245 120.635 56.415 120.805 ;
        RECT 56.705 120.635 56.875 120.805 ;
        RECT 57.165 120.635 57.335 120.805 ;
        RECT 57.625 120.635 57.795 120.805 ;
        RECT 58.085 120.635 58.255 120.805 ;
        RECT 58.545 120.635 58.715 120.805 ;
        RECT 59.005 120.635 59.175 120.805 ;
        RECT 59.465 120.635 59.635 120.805 ;
        RECT 59.925 120.635 60.095 120.805 ;
        RECT 60.385 120.635 60.555 120.805 ;
        RECT 60.845 120.635 61.015 120.805 ;
        RECT 61.305 120.635 61.475 120.805 ;
        RECT 61.765 120.635 61.935 120.805 ;
        RECT 62.225 120.635 62.395 120.805 ;
        RECT 62.685 120.635 62.855 120.805 ;
        RECT 63.145 120.635 63.315 120.805 ;
        RECT 63.605 120.635 63.775 120.805 ;
        RECT 64.065 120.635 64.235 120.805 ;
        RECT 64.525 120.635 64.695 120.805 ;
        RECT 64.985 120.635 65.155 120.805 ;
        RECT 65.445 120.635 65.615 120.805 ;
        RECT 65.905 120.635 66.075 120.805 ;
        RECT 66.365 120.635 66.535 120.805 ;
        RECT 66.825 120.635 66.995 120.805 ;
        RECT 67.285 120.635 67.455 120.805 ;
        RECT 67.745 120.635 67.915 120.805 ;
        RECT 68.205 120.635 68.375 120.805 ;
        RECT 68.665 120.635 68.835 120.805 ;
        RECT 69.125 120.635 69.295 120.805 ;
        RECT 69.585 120.635 69.755 120.805 ;
        RECT 70.045 120.635 70.215 120.805 ;
        RECT 70.505 120.635 70.675 120.805 ;
        RECT 70.965 120.635 71.135 120.805 ;
        RECT 71.425 120.635 71.595 120.805 ;
        RECT 71.885 120.635 72.055 120.805 ;
        RECT 72.345 120.635 72.515 120.805 ;
        RECT 72.805 120.635 72.975 120.805 ;
        RECT 73.265 120.635 73.435 120.805 ;
        RECT 73.725 120.635 73.895 120.805 ;
        RECT 74.185 120.635 74.355 120.805 ;
        RECT 74.645 120.635 74.815 120.805 ;
        RECT 75.105 120.635 75.275 120.805 ;
        RECT 75.565 120.635 75.735 120.805 ;
        RECT 76.025 120.635 76.195 120.805 ;
        RECT 76.485 120.635 76.655 120.805 ;
        RECT 76.945 120.635 77.115 120.805 ;
        RECT 77.405 120.635 77.575 120.805 ;
        RECT 77.865 120.635 78.035 120.805 ;
        RECT 78.325 120.635 78.495 120.805 ;
        RECT 78.785 120.635 78.955 120.805 ;
        RECT 79.245 120.635 79.415 120.805 ;
        RECT 79.705 120.635 79.875 120.805 ;
        RECT 80.165 120.635 80.335 120.805 ;
        RECT 80.625 120.635 80.795 120.805 ;
        RECT 81.085 120.635 81.255 120.805 ;
        RECT 81.545 120.635 81.715 120.805 ;
        RECT 82.005 120.635 82.175 120.805 ;
        RECT 82.465 120.635 82.635 120.805 ;
        RECT 82.925 120.635 83.095 120.805 ;
        RECT 83.385 120.635 83.555 120.805 ;
        RECT 83.845 120.635 84.015 120.805 ;
        RECT 84.305 120.635 84.475 120.805 ;
        RECT 84.765 120.635 84.935 120.805 ;
        RECT 85.225 120.635 85.395 120.805 ;
        RECT 85.685 120.635 85.855 120.805 ;
        RECT 86.145 120.635 86.315 120.805 ;
        RECT 86.605 120.635 86.775 120.805 ;
        RECT 87.065 120.635 87.235 120.805 ;
        RECT 87.525 120.635 87.695 120.805 ;
        RECT 87.985 120.635 88.155 120.805 ;
        RECT 88.445 120.635 88.615 120.805 ;
        RECT 88.905 120.635 89.075 120.805 ;
        RECT 89.365 120.635 89.535 120.805 ;
        RECT 89.825 120.635 89.995 120.805 ;
        RECT 90.285 120.635 90.455 120.805 ;
        RECT 90.745 120.635 90.915 120.805 ;
        RECT 91.205 120.635 91.375 120.805 ;
        RECT 91.665 120.635 91.835 120.805 ;
        RECT 92.125 120.635 92.295 120.805 ;
        RECT 92.585 120.635 92.755 120.805 ;
        RECT 93.045 120.635 93.215 120.805 ;
        RECT 93.505 120.635 93.675 120.805 ;
        RECT 93.965 120.635 94.135 120.805 ;
        RECT 94.425 120.635 94.595 120.805 ;
        RECT 94.885 120.635 95.055 120.805 ;
        RECT 95.345 120.635 95.515 120.805 ;
        RECT 95.805 120.635 95.975 120.805 ;
        RECT 96.265 120.635 96.435 120.805 ;
        RECT 96.725 120.635 96.895 120.805 ;
        RECT 97.185 120.635 97.355 120.805 ;
        RECT 97.645 120.635 97.815 120.805 ;
        RECT 98.105 120.635 98.275 120.805 ;
        RECT 98.565 120.635 98.735 120.805 ;
        RECT 99.025 120.635 99.195 120.805 ;
        RECT 99.485 120.635 99.655 120.805 ;
        RECT 99.945 120.635 100.115 120.805 ;
        RECT 100.405 120.635 100.575 120.805 ;
        RECT 100.865 120.635 101.035 120.805 ;
        RECT 101.325 120.635 101.495 120.805 ;
        RECT 101.785 120.635 101.955 120.805 ;
        RECT 102.245 120.635 102.415 120.805 ;
        RECT 102.705 120.635 102.875 120.805 ;
        RECT 103.165 120.635 103.335 120.805 ;
        RECT 103.625 120.635 103.795 120.805 ;
        RECT 104.085 120.635 104.255 120.805 ;
        RECT 104.545 120.635 104.715 120.805 ;
        RECT 105.005 120.635 105.175 120.805 ;
        RECT 105.465 120.635 105.635 120.805 ;
        RECT 105.925 120.635 106.095 120.805 ;
        RECT 106.385 120.635 106.555 120.805 ;
        RECT 106.845 120.635 107.015 120.805 ;
        RECT 107.305 120.635 107.475 120.805 ;
        RECT 107.765 120.635 107.935 120.805 ;
        RECT 108.225 120.635 108.395 120.805 ;
        RECT 108.685 120.635 108.855 120.805 ;
        RECT 109.145 120.635 109.315 120.805 ;
        RECT 109.605 120.635 109.775 120.805 ;
        RECT 110.065 120.635 110.235 120.805 ;
        RECT 110.525 120.635 110.695 120.805 ;
        RECT 110.985 120.635 111.155 120.805 ;
        RECT 111.445 120.635 111.615 120.805 ;
        RECT 111.905 120.635 112.075 120.805 ;
        RECT 112.365 120.635 112.535 120.805 ;
        RECT 112.825 120.635 112.995 120.805 ;
        RECT 113.285 120.635 113.455 120.805 ;
        RECT 113.745 120.635 113.915 120.805 ;
        RECT 114.205 120.635 114.375 120.805 ;
        RECT 114.665 120.635 114.835 120.805 ;
        RECT 115.125 120.635 115.295 120.805 ;
        RECT 115.585 120.635 115.755 120.805 ;
        RECT 116.045 120.635 116.215 120.805 ;
        RECT 116.505 120.635 116.675 120.805 ;
        RECT 116.965 120.635 117.135 120.805 ;
        RECT 117.425 120.635 117.595 120.805 ;
        RECT 117.885 120.635 118.055 120.805 ;
        RECT 118.345 120.635 118.515 120.805 ;
        RECT 118.805 120.635 118.975 120.805 ;
        RECT 119.265 120.635 119.435 120.805 ;
        RECT 119.725 120.635 119.895 120.805 ;
        RECT 120.185 120.635 120.355 120.805 ;
        RECT 120.645 120.635 120.815 120.805 ;
        RECT 121.105 120.635 121.275 120.805 ;
        RECT 121.565 120.635 121.735 120.805 ;
        RECT 122.025 120.635 122.195 120.805 ;
        RECT 122.485 120.635 122.655 120.805 ;
        RECT 122.945 120.635 123.115 120.805 ;
        RECT 123.405 120.635 123.575 120.805 ;
        RECT 123.865 120.635 124.035 120.805 ;
        RECT 124.325 120.635 124.495 120.805 ;
        RECT 124.785 120.635 124.955 120.805 ;
        RECT 125.245 120.635 125.415 120.805 ;
        RECT 125.705 120.635 125.875 120.805 ;
        RECT 126.165 120.635 126.335 120.805 ;
        RECT 126.625 120.635 126.795 120.805 ;
        RECT 127.085 120.635 127.255 120.805 ;
        RECT 127.545 120.635 127.715 120.805 ;
        RECT 128.005 120.635 128.175 120.805 ;
        RECT 128.465 120.635 128.635 120.805 ;
        RECT 128.925 120.635 129.095 120.805 ;
        RECT 129.385 120.635 129.555 120.805 ;
        RECT 129.845 120.635 130.015 120.805 ;
        RECT 130.305 120.635 130.475 120.805 ;
        RECT 130.765 120.635 130.935 120.805 ;
        RECT 131.225 120.635 131.395 120.805 ;
        RECT 131.685 120.635 131.855 120.805 ;
        RECT 132.145 120.635 132.315 120.805 ;
        RECT 132.605 120.635 132.775 120.805 ;
        RECT 133.065 120.635 133.235 120.805 ;
        RECT 133.525 120.635 133.695 120.805 ;
        RECT 133.985 120.635 134.155 120.805 ;
        RECT 45.665 115.195 45.835 115.365 ;
        RECT 46.125 115.195 46.295 115.365 ;
        RECT 46.585 115.195 46.755 115.365 ;
        RECT 47.045 115.195 47.215 115.365 ;
        RECT 47.505 115.195 47.675 115.365 ;
        RECT 47.965 115.195 48.135 115.365 ;
        RECT 48.425 115.195 48.595 115.365 ;
        RECT 48.885 115.195 49.055 115.365 ;
        RECT 49.345 115.195 49.515 115.365 ;
        RECT 49.805 115.195 49.975 115.365 ;
        RECT 50.265 115.195 50.435 115.365 ;
        RECT 50.725 115.195 50.895 115.365 ;
        RECT 51.185 115.195 51.355 115.365 ;
        RECT 51.645 115.195 51.815 115.365 ;
        RECT 52.105 115.195 52.275 115.365 ;
        RECT 52.565 115.195 52.735 115.365 ;
        RECT 53.025 115.195 53.195 115.365 ;
        RECT 53.485 115.195 53.655 115.365 ;
        RECT 53.945 115.195 54.115 115.365 ;
        RECT 54.405 115.195 54.575 115.365 ;
        RECT 54.865 115.195 55.035 115.365 ;
        RECT 55.325 115.195 55.495 115.365 ;
        RECT 55.785 115.195 55.955 115.365 ;
        RECT 56.245 115.195 56.415 115.365 ;
        RECT 56.705 115.195 56.875 115.365 ;
        RECT 57.165 115.195 57.335 115.365 ;
        RECT 57.625 115.195 57.795 115.365 ;
        RECT 58.085 115.195 58.255 115.365 ;
        RECT 58.545 115.195 58.715 115.365 ;
        RECT 59.005 115.195 59.175 115.365 ;
        RECT 59.465 115.195 59.635 115.365 ;
        RECT 59.925 115.195 60.095 115.365 ;
        RECT 60.385 115.195 60.555 115.365 ;
        RECT 60.845 115.195 61.015 115.365 ;
        RECT 61.305 115.195 61.475 115.365 ;
        RECT 61.765 115.195 61.935 115.365 ;
        RECT 62.225 115.195 62.395 115.365 ;
        RECT 62.685 115.195 62.855 115.365 ;
        RECT 63.145 115.195 63.315 115.365 ;
        RECT 63.605 115.195 63.775 115.365 ;
        RECT 64.065 115.195 64.235 115.365 ;
        RECT 64.525 115.195 64.695 115.365 ;
        RECT 64.985 115.195 65.155 115.365 ;
        RECT 65.445 115.195 65.615 115.365 ;
        RECT 65.905 115.195 66.075 115.365 ;
        RECT 66.365 115.195 66.535 115.365 ;
        RECT 66.825 115.195 66.995 115.365 ;
        RECT 67.285 115.195 67.455 115.365 ;
        RECT 67.745 115.195 67.915 115.365 ;
        RECT 68.205 115.195 68.375 115.365 ;
        RECT 68.665 115.195 68.835 115.365 ;
        RECT 69.125 115.195 69.295 115.365 ;
        RECT 69.585 115.195 69.755 115.365 ;
        RECT 70.045 115.195 70.215 115.365 ;
        RECT 70.505 115.195 70.675 115.365 ;
        RECT 70.965 115.195 71.135 115.365 ;
        RECT 71.425 115.195 71.595 115.365 ;
        RECT 71.885 115.195 72.055 115.365 ;
        RECT 72.345 115.195 72.515 115.365 ;
        RECT 72.805 115.195 72.975 115.365 ;
        RECT 73.265 115.195 73.435 115.365 ;
        RECT 73.725 115.195 73.895 115.365 ;
        RECT 74.185 115.195 74.355 115.365 ;
        RECT 74.645 115.195 74.815 115.365 ;
        RECT 75.105 115.195 75.275 115.365 ;
        RECT 75.565 115.195 75.735 115.365 ;
        RECT 76.025 115.195 76.195 115.365 ;
        RECT 76.485 115.195 76.655 115.365 ;
        RECT 76.945 115.195 77.115 115.365 ;
        RECT 77.405 115.195 77.575 115.365 ;
        RECT 77.865 115.195 78.035 115.365 ;
        RECT 78.325 115.195 78.495 115.365 ;
        RECT 78.785 115.195 78.955 115.365 ;
        RECT 79.245 115.195 79.415 115.365 ;
        RECT 79.705 115.195 79.875 115.365 ;
        RECT 80.165 115.195 80.335 115.365 ;
        RECT 80.625 115.195 80.795 115.365 ;
        RECT 81.085 115.195 81.255 115.365 ;
        RECT 81.545 115.195 81.715 115.365 ;
        RECT 82.005 115.195 82.175 115.365 ;
        RECT 82.465 115.195 82.635 115.365 ;
        RECT 82.925 115.195 83.095 115.365 ;
        RECT 83.385 115.195 83.555 115.365 ;
        RECT 83.845 115.195 84.015 115.365 ;
        RECT 84.305 115.195 84.475 115.365 ;
        RECT 84.765 115.195 84.935 115.365 ;
        RECT 85.225 115.195 85.395 115.365 ;
        RECT 85.685 115.195 85.855 115.365 ;
        RECT 86.145 115.195 86.315 115.365 ;
        RECT 86.605 115.195 86.775 115.365 ;
        RECT 87.065 115.195 87.235 115.365 ;
        RECT 87.525 115.195 87.695 115.365 ;
        RECT 87.985 115.195 88.155 115.365 ;
        RECT 88.445 115.195 88.615 115.365 ;
        RECT 88.905 115.195 89.075 115.365 ;
        RECT 89.365 115.195 89.535 115.365 ;
        RECT 89.825 115.195 89.995 115.365 ;
        RECT 90.285 115.195 90.455 115.365 ;
        RECT 90.745 115.195 90.915 115.365 ;
        RECT 91.205 115.195 91.375 115.365 ;
        RECT 91.665 115.195 91.835 115.365 ;
        RECT 92.125 115.195 92.295 115.365 ;
        RECT 92.585 115.195 92.755 115.365 ;
        RECT 93.045 115.195 93.215 115.365 ;
        RECT 93.505 115.195 93.675 115.365 ;
        RECT 93.965 115.195 94.135 115.365 ;
        RECT 94.425 115.195 94.595 115.365 ;
        RECT 94.885 115.195 95.055 115.365 ;
        RECT 95.345 115.195 95.515 115.365 ;
        RECT 95.805 115.195 95.975 115.365 ;
        RECT 96.265 115.195 96.435 115.365 ;
        RECT 96.725 115.195 96.895 115.365 ;
        RECT 97.185 115.195 97.355 115.365 ;
        RECT 97.645 115.195 97.815 115.365 ;
        RECT 98.105 115.195 98.275 115.365 ;
        RECT 98.565 115.195 98.735 115.365 ;
        RECT 99.025 115.195 99.195 115.365 ;
        RECT 99.485 115.195 99.655 115.365 ;
        RECT 99.945 115.195 100.115 115.365 ;
        RECT 100.405 115.195 100.575 115.365 ;
        RECT 100.865 115.195 101.035 115.365 ;
        RECT 101.325 115.195 101.495 115.365 ;
        RECT 101.785 115.195 101.955 115.365 ;
        RECT 102.245 115.195 102.415 115.365 ;
        RECT 102.705 115.195 102.875 115.365 ;
        RECT 103.165 115.195 103.335 115.365 ;
        RECT 103.625 115.195 103.795 115.365 ;
        RECT 104.085 115.195 104.255 115.365 ;
        RECT 104.545 115.195 104.715 115.365 ;
        RECT 105.005 115.195 105.175 115.365 ;
        RECT 105.465 115.195 105.635 115.365 ;
        RECT 105.925 115.195 106.095 115.365 ;
        RECT 106.385 115.195 106.555 115.365 ;
        RECT 106.845 115.195 107.015 115.365 ;
        RECT 107.305 115.195 107.475 115.365 ;
        RECT 107.765 115.195 107.935 115.365 ;
        RECT 108.225 115.195 108.395 115.365 ;
        RECT 108.685 115.195 108.855 115.365 ;
        RECT 109.145 115.195 109.315 115.365 ;
        RECT 109.605 115.195 109.775 115.365 ;
        RECT 110.065 115.195 110.235 115.365 ;
        RECT 110.525 115.195 110.695 115.365 ;
        RECT 110.985 115.195 111.155 115.365 ;
        RECT 111.445 115.195 111.615 115.365 ;
        RECT 111.905 115.195 112.075 115.365 ;
        RECT 112.365 115.195 112.535 115.365 ;
        RECT 112.825 115.195 112.995 115.365 ;
        RECT 113.285 115.195 113.455 115.365 ;
        RECT 113.745 115.195 113.915 115.365 ;
        RECT 114.205 115.195 114.375 115.365 ;
        RECT 114.665 115.195 114.835 115.365 ;
        RECT 115.125 115.195 115.295 115.365 ;
        RECT 115.585 115.195 115.755 115.365 ;
        RECT 116.045 115.195 116.215 115.365 ;
        RECT 116.505 115.195 116.675 115.365 ;
        RECT 116.965 115.195 117.135 115.365 ;
        RECT 117.425 115.195 117.595 115.365 ;
        RECT 117.885 115.195 118.055 115.365 ;
        RECT 118.345 115.195 118.515 115.365 ;
        RECT 118.805 115.195 118.975 115.365 ;
        RECT 119.265 115.195 119.435 115.365 ;
        RECT 119.725 115.195 119.895 115.365 ;
        RECT 120.185 115.195 120.355 115.365 ;
        RECT 120.645 115.195 120.815 115.365 ;
        RECT 121.105 115.195 121.275 115.365 ;
        RECT 121.565 115.195 121.735 115.365 ;
        RECT 122.025 115.195 122.195 115.365 ;
        RECT 122.485 115.195 122.655 115.365 ;
        RECT 122.945 115.195 123.115 115.365 ;
        RECT 123.405 115.195 123.575 115.365 ;
        RECT 123.865 115.195 124.035 115.365 ;
        RECT 124.325 115.195 124.495 115.365 ;
        RECT 124.785 115.195 124.955 115.365 ;
        RECT 125.245 115.195 125.415 115.365 ;
        RECT 125.705 115.195 125.875 115.365 ;
        RECT 126.165 115.195 126.335 115.365 ;
        RECT 126.625 115.195 126.795 115.365 ;
        RECT 127.085 115.195 127.255 115.365 ;
        RECT 127.545 115.195 127.715 115.365 ;
        RECT 128.005 115.195 128.175 115.365 ;
        RECT 128.465 115.195 128.635 115.365 ;
        RECT 128.925 115.195 129.095 115.365 ;
        RECT 129.385 115.195 129.555 115.365 ;
        RECT 129.845 115.195 130.015 115.365 ;
        RECT 130.305 115.195 130.475 115.365 ;
        RECT 130.765 115.195 130.935 115.365 ;
        RECT 131.225 115.195 131.395 115.365 ;
        RECT 131.685 115.195 131.855 115.365 ;
        RECT 132.145 115.195 132.315 115.365 ;
        RECT 132.605 115.195 132.775 115.365 ;
        RECT 133.065 115.195 133.235 115.365 ;
        RECT 133.525 115.195 133.695 115.365 ;
        RECT 133.985 115.195 134.155 115.365 ;
        RECT 45.665 109.755 45.835 109.925 ;
        RECT 46.125 109.755 46.295 109.925 ;
        RECT 46.585 109.755 46.755 109.925 ;
        RECT 47.045 109.755 47.215 109.925 ;
        RECT 47.505 109.755 47.675 109.925 ;
        RECT 47.965 109.755 48.135 109.925 ;
        RECT 48.425 109.755 48.595 109.925 ;
        RECT 48.885 109.755 49.055 109.925 ;
        RECT 49.345 109.755 49.515 109.925 ;
        RECT 49.805 109.755 49.975 109.925 ;
        RECT 50.265 109.755 50.435 109.925 ;
        RECT 50.725 109.755 50.895 109.925 ;
        RECT 51.185 109.755 51.355 109.925 ;
        RECT 51.645 109.755 51.815 109.925 ;
        RECT 52.105 109.755 52.275 109.925 ;
        RECT 52.565 109.755 52.735 109.925 ;
        RECT 53.025 109.755 53.195 109.925 ;
        RECT 53.485 109.755 53.655 109.925 ;
        RECT 53.945 109.755 54.115 109.925 ;
        RECT 54.405 109.755 54.575 109.925 ;
        RECT 54.865 109.755 55.035 109.925 ;
        RECT 55.325 109.755 55.495 109.925 ;
        RECT 55.785 109.755 55.955 109.925 ;
        RECT 56.245 109.755 56.415 109.925 ;
        RECT 56.705 109.755 56.875 109.925 ;
        RECT 57.165 109.755 57.335 109.925 ;
        RECT 57.625 109.755 57.795 109.925 ;
        RECT 58.085 109.755 58.255 109.925 ;
        RECT 58.545 109.755 58.715 109.925 ;
        RECT 59.005 109.755 59.175 109.925 ;
        RECT 59.465 109.755 59.635 109.925 ;
        RECT 59.925 109.755 60.095 109.925 ;
        RECT 60.385 109.755 60.555 109.925 ;
        RECT 60.845 109.755 61.015 109.925 ;
        RECT 61.305 109.755 61.475 109.925 ;
        RECT 61.765 109.755 61.935 109.925 ;
        RECT 62.225 109.755 62.395 109.925 ;
        RECT 62.685 109.755 62.855 109.925 ;
        RECT 63.145 109.755 63.315 109.925 ;
        RECT 63.605 109.755 63.775 109.925 ;
        RECT 64.065 109.755 64.235 109.925 ;
        RECT 64.525 109.755 64.695 109.925 ;
        RECT 64.985 109.755 65.155 109.925 ;
        RECT 65.445 109.755 65.615 109.925 ;
        RECT 65.905 109.755 66.075 109.925 ;
        RECT 66.365 109.755 66.535 109.925 ;
        RECT 66.825 109.755 66.995 109.925 ;
        RECT 67.285 109.755 67.455 109.925 ;
        RECT 67.745 109.755 67.915 109.925 ;
        RECT 68.205 109.755 68.375 109.925 ;
        RECT 68.665 109.755 68.835 109.925 ;
        RECT 69.125 109.755 69.295 109.925 ;
        RECT 69.585 109.755 69.755 109.925 ;
        RECT 70.045 109.755 70.215 109.925 ;
        RECT 70.505 109.755 70.675 109.925 ;
        RECT 70.965 109.755 71.135 109.925 ;
        RECT 71.425 109.755 71.595 109.925 ;
        RECT 71.885 109.755 72.055 109.925 ;
        RECT 72.345 109.755 72.515 109.925 ;
        RECT 72.805 109.755 72.975 109.925 ;
        RECT 73.265 109.755 73.435 109.925 ;
        RECT 73.725 109.755 73.895 109.925 ;
        RECT 74.185 109.755 74.355 109.925 ;
        RECT 74.645 109.755 74.815 109.925 ;
        RECT 75.105 109.755 75.275 109.925 ;
        RECT 75.565 109.755 75.735 109.925 ;
        RECT 76.025 109.755 76.195 109.925 ;
        RECT 76.485 109.755 76.655 109.925 ;
        RECT 76.945 109.755 77.115 109.925 ;
        RECT 77.405 109.755 77.575 109.925 ;
        RECT 77.865 109.755 78.035 109.925 ;
        RECT 78.325 109.755 78.495 109.925 ;
        RECT 78.785 109.755 78.955 109.925 ;
        RECT 79.245 109.755 79.415 109.925 ;
        RECT 79.705 109.755 79.875 109.925 ;
        RECT 80.165 109.755 80.335 109.925 ;
        RECT 80.625 109.755 80.795 109.925 ;
        RECT 81.085 109.755 81.255 109.925 ;
        RECT 81.545 109.755 81.715 109.925 ;
        RECT 82.005 109.755 82.175 109.925 ;
        RECT 82.465 109.755 82.635 109.925 ;
        RECT 82.925 109.755 83.095 109.925 ;
        RECT 83.385 109.755 83.555 109.925 ;
        RECT 83.845 109.755 84.015 109.925 ;
        RECT 84.305 109.755 84.475 109.925 ;
        RECT 84.765 109.755 84.935 109.925 ;
        RECT 85.225 109.755 85.395 109.925 ;
        RECT 85.685 109.755 85.855 109.925 ;
        RECT 86.145 109.755 86.315 109.925 ;
        RECT 86.605 109.755 86.775 109.925 ;
        RECT 87.065 109.755 87.235 109.925 ;
        RECT 87.525 109.755 87.695 109.925 ;
        RECT 87.985 109.755 88.155 109.925 ;
        RECT 88.445 109.755 88.615 109.925 ;
        RECT 88.905 109.755 89.075 109.925 ;
        RECT 89.365 109.755 89.535 109.925 ;
        RECT 89.825 109.755 89.995 109.925 ;
        RECT 90.285 109.755 90.455 109.925 ;
        RECT 90.745 109.755 90.915 109.925 ;
        RECT 91.205 109.755 91.375 109.925 ;
        RECT 91.665 109.755 91.835 109.925 ;
        RECT 92.125 109.755 92.295 109.925 ;
        RECT 92.585 109.755 92.755 109.925 ;
        RECT 93.045 109.755 93.215 109.925 ;
        RECT 93.505 109.755 93.675 109.925 ;
        RECT 93.965 109.755 94.135 109.925 ;
        RECT 94.425 109.755 94.595 109.925 ;
        RECT 94.885 109.755 95.055 109.925 ;
        RECT 95.345 109.755 95.515 109.925 ;
        RECT 95.805 109.755 95.975 109.925 ;
        RECT 96.265 109.755 96.435 109.925 ;
        RECT 96.725 109.755 96.895 109.925 ;
        RECT 97.185 109.755 97.355 109.925 ;
        RECT 97.645 109.755 97.815 109.925 ;
        RECT 98.105 109.755 98.275 109.925 ;
        RECT 98.565 109.755 98.735 109.925 ;
        RECT 99.025 109.755 99.195 109.925 ;
        RECT 99.485 109.755 99.655 109.925 ;
        RECT 99.945 109.755 100.115 109.925 ;
        RECT 100.405 109.755 100.575 109.925 ;
        RECT 100.865 109.755 101.035 109.925 ;
        RECT 101.325 109.755 101.495 109.925 ;
        RECT 101.785 109.755 101.955 109.925 ;
        RECT 102.245 109.755 102.415 109.925 ;
        RECT 102.705 109.755 102.875 109.925 ;
        RECT 103.165 109.755 103.335 109.925 ;
        RECT 103.625 109.755 103.795 109.925 ;
        RECT 104.085 109.755 104.255 109.925 ;
        RECT 104.545 109.755 104.715 109.925 ;
        RECT 105.005 109.755 105.175 109.925 ;
        RECT 105.465 109.755 105.635 109.925 ;
        RECT 105.925 109.755 106.095 109.925 ;
        RECT 106.385 109.755 106.555 109.925 ;
        RECT 106.845 109.755 107.015 109.925 ;
        RECT 107.305 109.755 107.475 109.925 ;
        RECT 107.765 109.755 107.935 109.925 ;
        RECT 108.225 109.755 108.395 109.925 ;
        RECT 108.685 109.755 108.855 109.925 ;
        RECT 109.145 109.755 109.315 109.925 ;
        RECT 109.605 109.755 109.775 109.925 ;
        RECT 110.065 109.755 110.235 109.925 ;
        RECT 110.525 109.755 110.695 109.925 ;
        RECT 110.985 109.755 111.155 109.925 ;
        RECT 111.445 109.755 111.615 109.925 ;
        RECT 111.905 109.755 112.075 109.925 ;
        RECT 112.365 109.755 112.535 109.925 ;
        RECT 112.825 109.755 112.995 109.925 ;
        RECT 113.285 109.755 113.455 109.925 ;
        RECT 113.745 109.755 113.915 109.925 ;
        RECT 114.205 109.755 114.375 109.925 ;
        RECT 114.665 109.755 114.835 109.925 ;
        RECT 115.125 109.755 115.295 109.925 ;
        RECT 115.585 109.755 115.755 109.925 ;
        RECT 116.045 109.755 116.215 109.925 ;
        RECT 116.505 109.755 116.675 109.925 ;
        RECT 116.965 109.755 117.135 109.925 ;
        RECT 117.425 109.755 117.595 109.925 ;
        RECT 117.885 109.755 118.055 109.925 ;
        RECT 118.345 109.755 118.515 109.925 ;
        RECT 118.805 109.755 118.975 109.925 ;
        RECT 119.265 109.755 119.435 109.925 ;
        RECT 119.725 109.755 119.895 109.925 ;
        RECT 120.185 109.755 120.355 109.925 ;
        RECT 120.645 109.755 120.815 109.925 ;
        RECT 121.105 109.755 121.275 109.925 ;
        RECT 121.565 109.755 121.735 109.925 ;
        RECT 122.025 109.755 122.195 109.925 ;
        RECT 122.485 109.755 122.655 109.925 ;
        RECT 122.945 109.755 123.115 109.925 ;
        RECT 123.405 109.755 123.575 109.925 ;
        RECT 123.865 109.755 124.035 109.925 ;
        RECT 124.325 109.755 124.495 109.925 ;
        RECT 124.785 109.755 124.955 109.925 ;
        RECT 125.245 109.755 125.415 109.925 ;
        RECT 125.705 109.755 125.875 109.925 ;
        RECT 126.165 109.755 126.335 109.925 ;
        RECT 126.625 109.755 126.795 109.925 ;
        RECT 127.085 109.755 127.255 109.925 ;
        RECT 127.545 109.755 127.715 109.925 ;
        RECT 128.005 109.755 128.175 109.925 ;
        RECT 128.465 109.755 128.635 109.925 ;
        RECT 128.925 109.755 129.095 109.925 ;
        RECT 129.385 109.755 129.555 109.925 ;
        RECT 129.845 109.755 130.015 109.925 ;
        RECT 130.305 109.755 130.475 109.925 ;
        RECT 130.765 109.755 130.935 109.925 ;
        RECT 131.225 109.755 131.395 109.925 ;
        RECT 131.685 109.755 131.855 109.925 ;
        RECT 132.145 109.755 132.315 109.925 ;
        RECT 132.605 109.755 132.775 109.925 ;
        RECT 133.065 109.755 133.235 109.925 ;
        RECT 133.525 109.755 133.695 109.925 ;
        RECT 133.985 109.755 134.155 109.925 ;
        RECT 45.665 104.315 45.835 104.485 ;
        RECT 46.125 104.315 46.295 104.485 ;
        RECT 46.585 104.315 46.755 104.485 ;
        RECT 47.045 104.315 47.215 104.485 ;
        RECT 47.505 104.315 47.675 104.485 ;
        RECT 47.965 104.315 48.135 104.485 ;
        RECT 48.425 104.315 48.595 104.485 ;
        RECT 48.885 104.315 49.055 104.485 ;
        RECT 49.345 104.315 49.515 104.485 ;
        RECT 49.805 104.315 49.975 104.485 ;
        RECT 50.265 104.315 50.435 104.485 ;
        RECT 50.725 104.315 50.895 104.485 ;
        RECT 51.185 104.315 51.355 104.485 ;
        RECT 51.645 104.315 51.815 104.485 ;
        RECT 52.105 104.315 52.275 104.485 ;
        RECT 52.565 104.315 52.735 104.485 ;
        RECT 53.025 104.315 53.195 104.485 ;
        RECT 53.485 104.315 53.655 104.485 ;
        RECT 53.945 104.315 54.115 104.485 ;
        RECT 54.405 104.315 54.575 104.485 ;
        RECT 54.865 104.315 55.035 104.485 ;
        RECT 55.325 104.315 55.495 104.485 ;
        RECT 55.785 104.315 55.955 104.485 ;
        RECT 56.245 104.315 56.415 104.485 ;
        RECT 56.705 104.315 56.875 104.485 ;
        RECT 57.165 104.315 57.335 104.485 ;
        RECT 57.625 104.315 57.795 104.485 ;
        RECT 58.085 104.315 58.255 104.485 ;
        RECT 58.545 104.315 58.715 104.485 ;
        RECT 59.005 104.315 59.175 104.485 ;
        RECT 59.465 104.315 59.635 104.485 ;
        RECT 59.925 104.315 60.095 104.485 ;
        RECT 60.385 104.315 60.555 104.485 ;
        RECT 60.845 104.315 61.015 104.485 ;
        RECT 61.305 104.315 61.475 104.485 ;
        RECT 61.765 104.315 61.935 104.485 ;
        RECT 62.225 104.315 62.395 104.485 ;
        RECT 62.685 104.315 62.855 104.485 ;
        RECT 63.145 104.315 63.315 104.485 ;
        RECT 63.605 104.315 63.775 104.485 ;
        RECT 64.065 104.315 64.235 104.485 ;
        RECT 64.525 104.315 64.695 104.485 ;
        RECT 64.985 104.315 65.155 104.485 ;
        RECT 65.445 104.315 65.615 104.485 ;
        RECT 65.905 104.315 66.075 104.485 ;
        RECT 66.365 104.315 66.535 104.485 ;
        RECT 66.825 104.315 66.995 104.485 ;
        RECT 67.285 104.315 67.455 104.485 ;
        RECT 67.745 104.315 67.915 104.485 ;
        RECT 68.205 104.315 68.375 104.485 ;
        RECT 68.665 104.315 68.835 104.485 ;
        RECT 69.125 104.315 69.295 104.485 ;
        RECT 69.585 104.315 69.755 104.485 ;
        RECT 70.045 104.315 70.215 104.485 ;
        RECT 70.505 104.315 70.675 104.485 ;
        RECT 70.965 104.315 71.135 104.485 ;
        RECT 71.425 104.315 71.595 104.485 ;
        RECT 71.885 104.315 72.055 104.485 ;
        RECT 72.345 104.315 72.515 104.485 ;
        RECT 72.805 104.315 72.975 104.485 ;
        RECT 73.265 104.315 73.435 104.485 ;
        RECT 73.725 104.315 73.895 104.485 ;
        RECT 74.185 104.315 74.355 104.485 ;
        RECT 74.645 104.315 74.815 104.485 ;
        RECT 75.105 104.315 75.275 104.485 ;
        RECT 75.565 104.315 75.735 104.485 ;
        RECT 76.025 104.315 76.195 104.485 ;
        RECT 76.485 104.315 76.655 104.485 ;
        RECT 76.945 104.315 77.115 104.485 ;
        RECT 77.405 104.315 77.575 104.485 ;
        RECT 77.865 104.315 78.035 104.485 ;
        RECT 78.325 104.315 78.495 104.485 ;
        RECT 78.785 104.315 78.955 104.485 ;
        RECT 79.245 104.315 79.415 104.485 ;
        RECT 79.705 104.315 79.875 104.485 ;
        RECT 80.165 104.315 80.335 104.485 ;
        RECT 80.625 104.315 80.795 104.485 ;
        RECT 81.085 104.315 81.255 104.485 ;
        RECT 81.545 104.315 81.715 104.485 ;
        RECT 82.005 104.315 82.175 104.485 ;
        RECT 82.465 104.315 82.635 104.485 ;
        RECT 82.925 104.315 83.095 104.485 ;
        RECT 83.385 104.315 83.555 104.485 ;
        RECT 83.845 104.315 84.015 104.485 ;
        RECT 84.305 104.315 84.475 104.485 ;
        RECT 84.765 104.315 84.935 104.485 ;
        RECT 85.225 104.315 85.395 104.485 ;
        RECT 85.685 104.315 85.855 104.485 ;
        RECT 86.145 104.315 86.315 104.485 ;
        RECT 86.605 104.315 86.775 104.485 ;
        RECT 87.065 104.315 87.235 104.485 ;
        RECT 87.525 104.315 87.695 104.485 ;
        RECT 87.985 104.315 88.155 104.485 ;
        RECT 88.445 104.315 88.615 104.485 ;
        RECT 88.905 104.315 89.075 104.485 ;
        RECT 89.365 104.315 89.535 104.485 ;
        RECT 89.825 104.315 89.995 104.485 ;
        RECT 90.285 104.315 90.455 104.485 ;
        RECT 90.745 104.315 90.915 104.485 ;
        RECT 91.205 104.315 91.375 104.485 ;
        RECT 91.665 104.315 91.835 104.485 ;
        RECT 92.125 104.315 92.295 104.485 ;
        RECT 92.585 104.315 92.755 104.485 ;
        RECT 93.045 104.315 93.215 104.485 ;
        RECT 93.505 104.315 93.675 104.485 ;
        RECT 93.965 104.315 94.135 104.485 ;
        RECT 94.425 104.315 94.595 104.485 ;
        RECT 94.885 104.315 95.055 104.485 ;
        RECT 95.345 104.315 95.515 104.485 ;
        RECT 95.805 104.315 95.975 104.485 ;
        RECT 96.265 104.315 96.435 104.485 ;
        RECT 96.725 104.315 96.895 104.485 ;
        RECT 97.185 104.315 97.355 104.485 ;
        RECT 97.645 104.315 97.815 104.485 ;
        RECT 98.105 104.315 98.275 104.485 ;
        RECT 98.565 104.315 98.735 104.485 ;
        RECT 99.025 104.315 99.195 104.485 ;
        RECT 99.485 104.315 99.655 104.485 ;
        RECT 99.945 104.315 100.115 104.485 ;
        RECT 100.405 104.315 100.575 104.485 ;
        RECT 100.865 104.315 101.035 104.485 ;
        RECT 101.325 104.315 101.495 104.485 ;
        RECT 101.785 104.315 101.955 104.485 ;
        RECT 102.245 104.315 102.415 104.485 ;
        RECT 102.705 104.315 102.875 104.485 ;
        RECT 103.165 104.315 103.335 104.485 ;
        RECT 103.625 104.315 103.795 104.485 ;
        RECT 104.085 104.315 104.255 104.485 ;
        RECT 104.545 104.315 104.715 104.485 ;
        RECT 105.005 104.315 105.175 104.485 ;
        RECT 105.465 104.315 105.635 104.485 ;
        RECT 105.925 104.315 106.095 104.485 ;
        RECT 106.385 104.315 106.555 104.485 ;
        RECT 106.845 104.315 107.015 104.485 ;
        RECT 107.305 104.315 107.475 104.485 ;
        RECT 107.765 104.315 107.935 104.485 ;
        RECT 108.225 104.315 108.395 104.485 ;
        RECT 108.685 104.315 108.855 104.485 ;
        RECT 109.145 104.315 109.315 104.485 ;
        RECT 109.605 104.315 109.775 104.485 ;
        RECT 110.065 104.315 110.235 104.485 ;
        RECT 110.525 104.315 110.695 104.485 ;
        RECT 110.985 104.315 111.155 104.485 ;
        RECT 111.445 104.315 111.615 104.485 ;
        RECT 111.905 104.315 112.075 104.485 ;
        RECT 112.365 104.315 112.535 104.485 ;
        RECT 112.825 104.315 112.995 104.485 ;
        RECT 113.285 104.315 113.455 104.485 ;
        RECT 113.745 104.315 113.915 104.485 ;
        RECT 114.205 104.315 114.375 104.485 ;
        RECT 114.665 104.315 114.835 104.485 ;
        RECT 115.125 104.315 115.295 104.485 ;
        RECT 115.585 104.315 115.755 104.485 ;
        RECT 116.045 104.315 116.215 104.485 ;
        RECT 116.505 104.315 116.675 104.485 ;
        RECT 116.965 104.315 117.135 104.485 ;
        RECT 117.425 104.315 117.595 104.485 ;
        RECT 117.885 104.315 118.055 104.485 ;
        RECT 118.345 104.315 118.515 104.485 ;
        RECT 118.805 104.315 118.975 104.485 ;
        RECT 119.265 104.315 119.435 104.485 ;
        RECT 119.725 104.315 119.895 104.485 ;
        RECT 120.185 104.315 120.355 104.485 ;
        RECT 120.645 104.315 120.815 104.485 ;
        RECT 121.105 104.315 121.275 104.485 ;
        RECT 121.565 104.315 121.735 104.485 ;
        RECT 122.025 104.315 122.195 104.485 ;
        RECT 122.485 104.315 122.655 104.485 ;
        RECT 122.945 104.315 123.115 104.485 ;
        RECT 123.405 104.315 123.575 104.485 ;
        RECT 123.865 104.315 124.035 104.485 ;
        RECT 124.325 104.315 124.495 104.485 ;
        RECT 124.785 104.315 124.955 104.485 ;
        RECT 125.245 104.315 125.415 104.485 ;
        RECT 125.705 104.315 125.875 104.485 ;
        RECT 126.165 104.315 126.335 104.485 ;
        RECT 126.625 104.315 126.795 104.485 ;
        RECT 127.085 104.315 127.255 104.485 ;
        RECT 127.545 104.315 127.715 104.485 ;
        RECT 128.005 104.315 128.175 104.485 ;
        RECT 128.465 104.315 128.635 104.485 ;
        RECT 128.925 104.315 129.095 104.485 ;
        RECT 129.385 104.315 129.555 104.485 ;
        RECT 129.845 104.315 130.015 104.485 ;
        RECT 130.305 104.315 130.475 104.485 ;
        RECT 130.765 104.315 130.935 104.485 ;
        RECT 131.225 104.315 131.395 104.485 ;
        RECT 131.685 104.315 131.855 104.485 ;
        RECT 132.145 104.315 132.315 104.485 ;
        RECT 132.605 104.315 132.775 104.485 ;
        RECT 133.065 104.315 133.235 104.485 ;
        RECT 133.525 104.315 133.695 104.485 ;
        RECT 133.985 104.315 134.155 104.485 ;
        RECT 45.665 98.875 45.835 99.045 ;
        RECT 46.125 98.875 46.295 99.045 ;
        RECT 46.585 98.875 46.755 99.045 ;
        RECT 47.045 98.875 47.215 99.045 ;
        RECT 47.505 98.875 47.675 99.045 ;
        RECT 47.965 98.875 48.135 99.045 ;
        RECT 48.425 98.875 48.595 99.045 ;
        RECT 48.885 98.875 49.055 99.045 ;
        RECT 49.345 98.875 49.515 99.045 ;
        RECT 49.805 98.875 49.975 99.045 ;
        RECT 50.265 98.875 50.435 99.045 ;
        RECT 50.725 98.875 50.895 99.045 ;
        RECT 51.185 98.875 51.355 99.045 ;
        RECT 51.645 98.875 51.815 99.045 ;
        RECT 52.105 98.875 52.275 99.045 ;
        RECT 52.565 98.875 52.735 99.045 ;
        RECT 53.025 98.875 53.195 99.045 ;
        RECT 53.485 98.875 53.655 99.045 ;
        RECT 53.945 98.875 54.115 99.045 ;
        RECT 54.405 98.875 54.575 99.045 ;
        RECT 54.865 98.875 55.035 99.045 ;
        RECT 55.325 98.875 55.495 99.045 ;
        RECT 55.785 98.875 55.955 99.045 ;
        RECT 56.245 98.875 56.415 99.045 ;
        RECT 56.705 98.875 56.875 99.045 ;
        RECT 57.165 98.875 57.335 99.045 ;
        RECT 57.625 98.875 57.795 99.045 ;
        RECT 58.085 98.875 58.255 99.045 ;
        RECT 58.545 98.875 58.715 99.045 ;
        RECT 59.005 98.875 59.175 99.045 ;
        RECT 59.465 98.875 59.635 99.045 ;
        RECT 59.925 98.875 60.095 99.045 ;
        RECT 60.385 98.875 60.555 99.045 ;
        RECT 60.845 98.875 61.015 99.045 ;
        RECT 61.305 98.875 61.475 99.045 ;
        RECT 61.765 98.875 61.935 99.045 ;
        RECT 62.225 98.875 62.395 99.045 ;
        RECT 62.685 98.875 62.855 99.045 ;
        RECT 63.145 98.875 63.315 99.045 ;
        RECT 63.605 98.875 63.775 99.045 ;
        RECT 64.065 98.875 64.235 99.045 ;
        RECT 64.525 98.875 64.695 99.045 ;
        RECT 64.985 98.875 65.155 99.045 ;
        RECT 65.445 98.875 65.615 99.045 ;
        RECT 65.905 98.875 66.075 99.045 ;
        RECT 66.365 98.875 66.535 99.045 ;
        RECT 66.825 98.875 66.995 99.045 ;
        RECT 67.285 98.875 67.455 99.045 ;
        RECT 67.745 98.875 67.915 99.045 ;
        RECT 68.205 98.875 68.375 99.045 ;
        RECT 68.665 98.875 68.835 99.045 ;
        RECT 69.125 98.875 69.295 99.045 ;
        RECT 69.585 98.875 69.755 99.045 ;
        RECT 70.045 98.875 70.215 99.045 ;
        RECT 70.505 98.875 70.675 99.045 ;
        RECT 70.965 98.875 71.135 99.045 ;
        RECT 71.425 98.875 71.595 99.045 ;
        RECT 71.885 98.875 72.055 99.045 ;
        RECT 72.345 98.875 72.515 99.045 ;
        RECT 72.805 98.875 72.975 99.045 ;
        RECT 73.265 98.875 73.435 99.045 ;
        RECT 73.725 98.875 73.895 99.045 ;
        RECT 74.185 98.875 74.355 99.045 ;
        RECT 74.645 98.875 74.815 99.045 ;
        RECT 75.105 98.875 75.275 99.045 ;
        RECT 75.565 98.875 75.735 99.045 ;
        RECT 76.025 98.875 76.195 99.045 ;
        RECT 76.485 98.875 76.655 99.045 ;
        RECT 76.945 98.875 77.115 99.045 ;
        RECT 77.405 98.875 77.575 99.045 ;
        RECT 77.865 98.875 78.035 99.045 ;
        RECT 78.325 98.875 78.495 99.045 ;
        RECT 78.785 98.875 78.955 99.045 ;
        RECT 79.245 98.875 79.415 99.045 ;
        RECT 79.705 98.875 79.875 99.045 ;
        RECT 80.165 98.875 80.335 99.045 ;
        RECT 80.625 98.875 80.795 99.045 ;
        RECT 81.085 98.875 81.255 99.045 ;
        RECT 81.545 98.875 81.715 99.045 ;
        RECT 82.005 98.875 82.175 99.045 ;
        RECT 82.465 98.875 82.635 99.045 ;
        RECT 82.925 98.875 83.095 99.045 ;
        RECT 83.385 98.875 83.555 99.045 ;
        RECT 83.845 98.875 84.015 99.045 ;
        RECT 84.305 98.875 84.475 99.045 ;
        RECT 84.765 98.875 84.935 99.045 ;
        RECT 85.225 98.875 85.395 99.045 ;
        RECT 85.685 98.875 85.855 99.045 ;
        RECT 86.145 98.875 86.315 99.045 ;
        RECT 86.605 98.875 86.775 99.045 ;
        RECT 87.065 98.875 87.235 99.045 ;
        RECT 87.525 98.875 87.695 99.045 ;
        RECT 87.985 98.875 88.155 99.045 ;
        RECT 88.445 98.875 88.615 99.045 ;
        RECT 88.905 98.875 89.075 99.045 ;
        RECT 89.365 98.875 89.535 99.045 ;
        RECT 89.825 98.875 89.995 99.045 ;
        RECT 90.285 98.875 90.455 99.045 ;
        RECT 90.745 98.875 90.915 99.045 ;
        RECT 91.205 98.875 91.375 99.045 ;
        RECT 91.665 98.875 91.835 99.045 ;
        RECT 92.125 98.875 92.295 99.045 ;
        RECT 92.585 98.875 92.755 99.045 ;
        RECT 93.045 98.875 93.215 99.045 ;
        RECT 93.505 98.875 93.675 99.045 ;
        RECT 93.965 98.875 94.135 99.045 ;
        RECT 94.425 98.875 94.595 99.045 ;
        RECT 94.885 98.875 95.055 99.045 ;
        RECT 95.345 98.875 95.515 99.045 ;
        RECT 95.805 98.875 95.975 99.045 ;
        RECT 96.265 98.875 96.435 99.045 ;
        RECT 96.725 98.875 96.895 99.045 ;
        RECT 97.185 98.875 97.355 99.045 ;
        RECT 97.645 98.875 97.815 99.045 ;
        RECT 98.105 98.875 98.275 99.045 ;
        RECT 98.565 98.875 98.735 99.045 ;
        RECT 99.025 98.875 99.195 99.045 ;
        RECT 99.485 98.875 99.655 99.045 ;
        RECT 99.945 98.875 100.115 99.045 ;
        RECT 100.405 98.875 100.575 99.045 ;
        RECT 100.865 98.875 101.035 99.045 ;
        RECT 101.325 98.875 101.495 99.045 ;
        RECT 101.785 98.875 101.955 99.045 ;
        RECT 102.245 98.875 102.415 99.045 ;
        RECT 102.705 98.875 102.875 99.045 ;
        RECT 103.165 98.875 103.335 99.045 ;
        RECT 103.625 98.875 103.795 99.045 ;
        RECT 104.085 98.875 104.255 99.045 ;
        RECT 104.545 98.875 104.715 99.045 ;
        RECT 105.005 98.875 105.175 99.045 ;
        RECT 105.465 98.875 105.635 99.045 ;
        RECT 105.925 98.875 106.095 99.045 ;
        RECT 106.385 98.875 106.555 99.045 ;
        RECT 106.845 98.875 107.015 99.045 ;
        RECT 107.305 98.875 107.475 99.045 ;
        RECT 107.765 98.875 107.935 99.045 ;
        RECT 108.225 98.875 108.395 99.045 ;
        RECT 108.685 98.875 108.855 99.045 ;
        RECT 109.145 98.875 109.315 99.045 ;
        RECT 109.605 98.875 109.775 99.045 ;
        RECT 110.065 98.875 110.235 99.045 ;
        RECT 110.525 98.875 110.695 99.045 ;
        RECT 110.985 98.875 111.155 99.045 ;
        RECT 111.445 98.875 111.615 99.045 ;
        RECT 111.905 98.875 112.075 99.045 ;
        RECT 112.365 98.875 112.535 99.045 ;
        RECT 112.825 98.875 112.995 99.045 ;
        RECT 113.285 98.875 113.455 99.045 ;
        RECT 113.745 98.875 113.915 99.045 ;
        RECT 114.205 98.875 114.375 99.045 ;
        RECT 114.665 98.875 114.835 99.045 ;
        RECT 115.125 98.875 115.295 99.045 ;
        RECT 115.585 98.875 115.755 99.045 ;
        RECT 116.045 98.875 116.215 99.045 ;
        RECT 116.505 98.875 116.675 99.045 ;
        RECT 116.965 98.875 117.135 99.045 ;
        RECT 117.425 98.875 117.595 99.045 ;
        RECT 117.885 98.875 118.055 99.045 ;
        RECT 118.345 98.875 118.515 99.045 ;
        RECT 118.805 98.875 118.975 99.045 ;
        RECT 119.265 98.875 119.435 99.045 ;
        RECT 119.725 98.875 119.895 99.045 ;
        RECT 120.185 98.875 120.355 99.045 ;
        RECT 120.645 98.875 120.815 99.045 ;
        RECT 121.105 98.875 121.275 99.045 ;
        RECT 121.565 98.875 121.735 99.045 ;
        RECT 122.025 98.875 122.195 99.045 ;
        RECT 122.485 98.875 122.655 99.045 ;
        RECT 122.945 98.875 123.115 99.045 ;
        RECT 123.405 98.875 123.575 99.045 ;
        RECT 123.865 98.875 124.035 99.045 ;
        RECT 124.325 98.875 124.495 99.045 ;
        RECT 124.785 98.875 124.955 99.045 ;
        RECT 125.245 98.875 125.415 99.045 ;
        RECT 125.705 98.875 125.875 99.045 ;
        RECT 126.165 98.875 126.335 99.045 ;
        RECT 126.625 98.875 126.795 99.045 ;
        RECT 127.085 98.875 127.255 99.045 ;
        RECT 127.545 98.875 127.715 99.045 ;
        RECT 128.005 98.875 128.175 99.045 ;
        RECT 128.465 98.875 128.635 99.045 ;
        RECT 128.925 98.875 129.095 99.045 ;
        RECT 129.385 98.875 129.555 99.045 ;
        RECT 129.845 98.875 130.015 99.045 ;
        RECT 130.305 98.875 130.475 99.045 ;
        RECT 130.765 98.875 130.935 99.045 ;
        RECT 131.225 98.875 131.395 99.045 ;
        RECT 131.685 98.875 131.855 99.045 ;
        RECT 132.145 98.875 132.315 99.045 ;
        RECT 132.605 98.875 132.775 99.045 ;
        RECT 133.065 98.875 133.235 99.045 ;
        RECT 133.525 98.875 133.695 99.045 ;
        RECT 133.985 98.875 134.155 99.045 ;
        RECT 45.665 93.435 45.835 93.605 ;
        RECT 46.125 93.435 46.295 93.605 ;
        RECT 46.585 93.435 46.755 93.605 ;
        RECT 47.045 93.435 47.215 93.605 ;
        RECT 47.505 93.435 47.675 93.605 ;
        RECT 47.965 93.435 48.135 93.605 ;
        RECT 48.425 93.435 48.595 93.605 ;
        RECT 48.885 93.435 49.055 93.605 ;
        RECT 49.345 93.435 49.515 93.605 ;
        RECT 49.805 93.435 49.975 93.605 ;
        RECT 50.265 93.435 50.435 93.605 ;
        RECT 50.725 93.435 50.895 93.605 ;
        RECT 51.185 93.435 51.355 93.605 ;
        RECT 51.645 93.435 51.815 93.605 ;
        RECT 52.105 93.435 52.275 93.605 ;
        RECT 52.565 93.435 52.735 93.605 ;
        RECT 53.025 93.435 53.195 93.605 ;
        RECT 53.485 93.435 53.655 93.605 ;
        RECT 53.945 93.435 54.115 93.605 ;
        RECT 54.405 93.435 54.575 93.605 ;
        RECT 54.865 93.435 55.035 93.605 ;
        RECT 55.325 93.435 55.495 93.605 ;
        RECT 55.785 93.435 55.955 93.605 ;
        RECT 56.245 93.435 56.415 93.605 ;
        RECT 56.705 93.435 56.875 93.605 ;
        RECT 57.165 93.435 57.335 93.605 ;
        RECT 57.625 93.435 57.795 93.605 ;
        RECT 58.085 93.435 58.255 93.605 ;
        RECT 58.545 93.435 58.715 93.605 ;
        RECT 59.005 93.435 59.175 93.605 ;
        RECT 59.465 93.435 59.635 93.605 ;
        RECT 59.925 93.435 60.095 93.605 ;
        RECT 60.385 93.435 60.555 93.605 ;
        RECT 60.845 93.435 61.015 93.605 ;
        RECT 61.305 93.435 61.475 93.605 ;
        RECT 61.765 93.435 61.935 93.605 ;
        RECT 62.225 93.435 62.395 93.605 ;
        RECT 62.685 93.435 62.855 93.605 ;
        RECT 63.145 93.435 63.315 93.605 ;
        RECT 63.605 93.435 63.775 93.605 ;
        RECT 64.065 93.435 64.235 93.605 ;
        RECT 64.525 93.435 64.695 93.605 ;
        RECT 64.985 93.435 65.155 93.605 ;
        RECT 65.445 93.435 65.615 93.605 ;
        RECT 65.905 93.435 66.075 93.605 ;
        RECT 66.365 93.435 66.535 93.605 ;
        RECT 66.825 93.435 66.995 93.605 ;
        RECT 67.285 93.435 67.455 93.605 ;
        RECT 67.745 93.435 67.915 93.605 ;
        RECT 68.205 93.435 68.375 93.605 ;
        RECT 68.665 93.435 68.835 93.605 ;
        RECT 69.125 93.435 69.295 93.605 ;
        RECT 69.585 93.435 69.755 93.605 ;
        RECT 70.045 93.435 70.215 93.605 ;
        RECT 70.505 93.435 70.675 93.605 ;
        RECT 70.965 93.435 71.135 93.605 ;
        RECT 71.425 93.435 71.595 93.605 ;
        RECT 71.885 93.435 72.055 93.605 ;
        RECT 72.345 93.435 72.515 93.605 ;
        RECT 72.805 93.435 72.975 93.605 ;
        RECT 73.265 93.435 73.435 93.605 ;
        RECT 73.725 93.435 73.895 93.605 ;
        RECT 74.185 93.435 74.355 93.605 ;
        RECT 74.645 93.435 74.815 93.605 ;
        RECT 75.105 93.435 75.275 93.605 ;
        RECT 75.565 93.435 75.735 93.605 ;
        RECT 76.025 93.435 76.195 93.605 ;
        RECT 76.485 93.435 76.655 93.605 ;
        RECT 76.945 93.435 77.115 93.605 ;
        RECT 77.405 93.435 77.575 93.605 ;
        RECT 77.865 93.435 78.035 93.605 ;
        RECT 78.325 93.435 78.495 93.605 ;
        RECT 78.785 93.435 78.955 93.605 ;
        RECT 79.245 93.435 79.415 93.605 ;
        RECT 79.705 93.435 79.875 93.605 ;
        RECT 80.165 93.435 80.335 93.605 ;
        RECT 80.625 93.435 80.795 93.605 ;
        RECT 81.085 93.435 81.255 93.605 ;
        RECT 81.545 93.435 81.715 93.605 ;
        RECT 82.005 93.435 82.175 93.605 ;
        RECT 82.465 93.435 82.635 93.605 ;
        RECT 82.925 93.435 83.095 93.605 ;
        RECT 83.385 93.435 83.555 93.605 ;
        RECT 83.845 93.435 84.015 93.605 ;
        RECT 84.305 93.435 84.475 93.605 ;
        RECT 84.765 93.435 84.935 93.605 ;
        RECT 85.225 93.435 85.395 93.605 ;
        RECT 85.685 93.435 85.855 93.605 ;
        RECT 86.145 93.435 86.315 93.605 ;
        RECT 86.605 93.435 86.775 93.605 ;
        RECT 87.065 93.435 87.235 93.605 ;
        RECT 87.525 93.435 87.695 93.605 ;
        RECT 87.985 93.435 88.155 93.605 ;
        RECT 88.445 93.435 88.615 93.605 ;
        RECT 88.905 93.435 89.075 93.605 ;
        RECT 89.365 93.435 89.535 93.605 ;
        RECT 89.825 93.435 89.995 93.605 ;
        RECT 90.285 93.435 90.455 93.605 ;
        RECT 90.745 93.435 90.915 93.605 ;
        RECT 91.205 93.435 91.375 93.605 ;
        RECT 91.665 93.435 91.835 93.605 ;
        RECT 92.125 93.435 92.295 93.605 ;
        RECT 92.585 93.435 92.755 93.605 ;
        RECT 93.045 93.435 93.215 93.605 ;
        RECT 93.505 93.435 93.675 93.605 ;
        RECT 93.965 93.435 94.135 93.605 ;
        RECT 94.425 93.435 94.595 93.605 ;
        RECT 94.885 93.435 95.055 93.605 ;
        RECT 95.345 93.435 95.515 93.605 ;
        RECT 95.805 93.435 95.975 93.605 ;
        RECT 96.265 93.435 96.435 93.605 ;
        RECT 96.725 93.435 96.895 93.605 ;
        RECT 97.185 93.435 97.355 93.605 ;
        RECT 97.645 93.435 97.815 93.605 ;
        RECT 98.105 93.435 98.275 93.605 ;
        RECT 98.565 93.435 98.735 93.605 ;
        RECT 99.025 93.435 99.195 93.605 ;
        RECT 99.485 93.435 99.655 93.605 ;
        RECT 99.945 93.435 100.115 93.605 ;
        RECT 100.405 93.435 100.575 93.605 ;
        RECT 100.865 93.435 101.035 93.605 ;
        RECT 101.325 93.435 101.495 93.605 ;
        RECT 101.785 93.435 101.955 93.605 ;
        RECT 102.245 93.435 102.415 93.605 ;
        RECT 102.705 93.435 102.875 93.605 ;
        RECT 103.165 93.435 103.335 93.605 ;
        RECT 103.625 93.435 103.795 93.605 ;
        RECT 104.085 93.435 104.255 93.605 ;
        RECT 104.545 93.435 104.715 93.605 ;
        RECT 105.005 93.435 105.175 93.605 ;
        RECT 105.465 93.435 105.635 93.605 ;
        RECT 105.925 93.435 106.095 93.605 ;
        RECT 106.385 93.435 106.555 93.605 ;
        RECT 106.845 93.435 107.015 93.605 ;
        RECT 107.305 93.435 107.475 93.605 ;
        RECT 107.765 93.435 107.935 93.605 ;
        RECT 108.225 93.435 108.395 93.605 ;
        RECT 108.685 93.435 108.855 93.605 ;
        RECT 109.145 93.435 109.315 93.605 ;
        RECT 109.605 93.435 109.775 93.605 ;
        RECT 110.065 93.435 110.235 93.605 ;
        RECT 110.525 93.435 110.695 93.605 ;
        RECT 110.985 93.435 111.155 93.605 ;
        RECT 111.445 93.435 111.615 93.605 ;
        RECT 111.905 93.435 112.075 93.605 ;
        RECT 112.365 93.435 112.535 93.605 ;
        RECT 112.825 93.435 112.995 93.605 ;
        RECT 113.285 93.435 113.455 93.605 ;
        RECT 113.745 93.435 113.915 93.605 ;
        RECT 114.205 93.435 114.375 93.605 ;
        RECT 114.665 93.435 114.835 93.605 ;
        RECT 115.125 93.435 115.295 93.605 ;
        RECT 115.585 93.435 115.755 93.605 ;
        RECT 116.045 93.435 116.215 93.605 ;
        RECT 116.505 93.435 116.675 93.605 ;
        RECT 116.965 93.435 117.135 93.605 ;
        RECT 117.425 93.435 117.595 93.605 ;
        RECT 117.885 93.435 118.055 93.605 ;
        RECT 118.345 93.435 118.515 93.605 ;
        RECT 118.805 93.435 118.975 93.605 ;
        RECT 119.265 93.435 119.435 93.605 ;
        RECT 119.725 93.435 119.895 93.605 ;
        RECT 120.185 93.435 120.355 93.605 ;
        RECT 120.645 93.435 120.815 93.605 ;
        RECT 121.105 93.435 121.275 93.605 ;
        RECT 121.565 93.435 121.735 93.605 ;
        RECT 122.025 93.435 122.195 93.605 ;
        RECT 122.485 93.435 122.655 93.605 ;
        RECT 122.945 93.435 123.115 93.605 ;
        RECT 123.405 93.435 123.575 93.605 ;
        RECT 123.865 93.435 124.035 93.605 ;
        RECT 124.325 93.435 124.495 93.605 ;
        RECT 124.785 93.435 124.955 93.605 ;
        RECT 125.245 93.435 125.415 93.605 ;
        RECT 125.705 93.435 125.875 93.605 ;
        RECT 126.165 93.435 126.335 93.605 ;
        RECT 126.625 93.435 126.795 93.605 ;
        RECT 127.085 93.435 127.255 93.605 ;
        RECT 127.545 93.435 127.715 93.605 ;
        RECT 128.005 93.435 128.175 93.605 ;
        RECT 128.465 93.435 128.635 93.605 ;
        RECT 128.925 93.435 129.095 93.605 ;
        RECT 129.385 93.435 129.555 93.605 ;
        RECT 129.845 93.435 130.015 93.605 ;
        RECT 130.305 93.435 130.475 93.605 ;
        RECT 130.765 93.435 130.935 93.605 ;
        RECT 131.225 93.435 131.395 93.605 ;
        RECT 131.685 93.435 131.855 93.605 ;
        RECT 132.145 93.435 132.315 93.605 ;
        RECT 132.605 93.435 132.775 93.605 ;
        RECT 133.065 93.435 133.235 93.605 ;
        RECT 133.525 93.435 133.695 93.605 ;
        RECT 133.985 93.435 134.155 93.605 ;
        RECT 45.665 87.995 45.835 88.165 ;
        RECT 46.125 87.995 46.295 88.165 ;
        RECT 46.585 87.995 46.755 88.165 ;
        RECT 47.045 87.995 47.215 88.165 ;
        RECT 47.505 87.995 47.675 88.165 ;
        RECT 47.965 87.995 48.135 88.165 ;
        RECT 48.425 87.995 48.595 88.165 ;
        RECT 48.885 87.995 49.055 88.165 ;
        RECT 49.345 87.995 49.515 88.165 ;
        RECT 49.805 87.995 49.975 88.165 ;
        RECT 50.265 87.995 50.435 88.165 ;
        RECT 50.725 87.995 50.895 88.165 ;
        RECT 51.185 87.995 51.355 88.165 ;
        RECT 51.645 87.995 51.815 88.165 ;
        RECT 52.105 87.995 52.275 88.165 ;
        RECT 52.565 87.995 52.735 88.165 ;
        RECT 53.025 87.995 53.195 88.165 ;
        RECT 53.485 87.995 53.655 88.165 ;
        RECT 53.945 87.995 54.115 88.165 ;
        RECT 54.405 87.995 54.575 88.165 ;
        RECT 54.865 87.995 55.035 88.165 ;
        RECT 55.325 87.995 55.495 88.165 ;
        RECT 55.785 87.995 55.955 88.165 ;
        RECT 56.245 87.995 56.415 88.165 ;
        RECT 56.705 87.995 56.875 88.165 ;
        RECT 57.165 87.995 57.335 88.165 ;
        RECT 57.625 87.995 57.795 88.165 ;
        RECT 58.085 87.995 58.255 88.165 ;
        RECT 58.545 87.995 58.715 88.165 ;
        RECT 59.005 87.995 59.175 88.165 ;
        RECT 59.465 87.995 59.635 88.165 ;
        RECT 59.925 87.995 60.095 88.165 ;
        RECT 60.385 87.995 60.555 88.165 ;
        RECT 60.845 87.995 61.015 88.165 ;
        RECT 61.305 87.995 61.475 88.165 ;
        RECT 61.765 87.995 61.935 88.165 ;
        RECT 62.225 87.995 62.395 88.165 ;
        RECT 62.685 87.995 62.855 88.165 ;
        RECT 63.145 87.995 63.315 88.165 ;
        RECT 63.605 87.995 63.775 88.165 ;
        RECT 64.065 87.995 64.235 88.165 ;
        RECT 64.525 87.995 64.695 88.165 ;
        RECT 64.985 87.995 65.155 88.165 ;
        RECT 65.445 87.995 65.615 88.165 ;
        RECT 65.905 87.995 66.075 88.165 ;
        RECT 66.365 87.995 66.535 88.165 ;
        RECT 66.825 87.995 66.995 88.165 ;
        RECT 67.285 87.995 67.455 88.165 ;
        RECT 67.745 87.995 67.915 88.165 ;
        RECT 68.205 87.995 68.375 88.165 ;
        RECT 68.665 87.995 68.835 88.165 ;
        RECT 69.125 87.995 69.295 88.165 ;
        RECT 69.585 87.995 69.755 88.165 ;
        RECT 70.045 87.995 70.215 88.165 ;
        RECT 70.505 87.995 70.675 88.165 ;
        RECT 70.965 87.995 71.135 88.165 ;
        RECT 71.425 87.995 71.595 88.165 ;
        RECT 71.885 87.995 72.055 88.165 ;
        RECT 72.345 87.995 72.515 88.165 ;
        RECT 72.805 87.995 72.975 88.165 ;
        RECT 73.265 87.995 73.435 88.165 ;
        RECT 73.725 87.995 73.895 88.165 ;
        RECT 74.185 87.995 74.355 88.165 ;
        RECT 74.645 87.995 74.815 88.165 ;
        RECT 75.105 87.995 75.275 88.165 ;
        RECT 75.565 87.995 75.735 88.165 ;
        RECT 76.025 87.995 76.195 88.165 ;
        RECT 76.485 87.995 76.655 88.165 ;
        RECT 76.945 87.995 77.115 88.165 ;
        RECT 77.405 87.995 77.575 88.165 ;
        RECT 77.865 87.995 78.035 88.165 ;
        RECT 78.325 87.995 78.495 88.165 ;
        RECT 78.785 87.995 78.955 88.165 ;
        RECT 79.245 87.995 79.415 88.165 ;
        RECT 79.705 87.995 79.875 88.165 ;
        RECT 80.165 87.995 80.335 88.165 ;
        RECT 80.625 87.995 80.795 88.165 ;
        RECT 81.085 87.995 81.255 88.165 ;
        RECT 81.545 87.995 81.715 88.165 ;
        RECT 82.005 87.995 82.175 88.165 ;
        RECT 82.465 87.995 82.635 88.165 ;
        RECT 82.925 87.995 83.095 88.165 ;
        RECT 83.385 87.995 83.555 88.165 ;
        RECT 83.845 87.995 84.015 88.165 ;
        RECT 84.305 87.995 84.475 88.165 ;
        RECT 84.765 87.995 84.935 88.165 ;
        RECT 85.225 87.995 85.395 88.165 ;
        RECT 85.685 87.995 85.855 88.165 ;
        RECT 86.145 87.995 86.315 88.165 ;
        RECT 86.605 87.995 86.775 88.165 ;
        RECT 87.065 87.995 87.235 88.165 ;
        RECT 87.525 87.995 87.695 88.165 ;
        RECT 87.985 87.995 88.155 88.165 ;
        RECT 88.445 87.995 88.615 88.165 ;
        RECT 88.905 87.995 89.075 88.165 ;
        RECT 89.365 87.995 89.535 88.165 ;
        RECT 89.825 87.995 89.995 88.165 ;
        RECT 90.285 87.995 90.455 88.165 ;
        RECT 90.745 87.995 90.915 88.165 ;
        RECT 91.205 87.995 91.375 88.165 ;
        RECT 91.665 87.995 91.835 88.165 ;
        RECT 92.125 87.995 92.295 88.165 ;
        RECT 92.585 87.995 92.755 88.165 ;
        RECT 93.045 87.995 93.215 88.165 ;
        RECT 93.505 87.995 93.675 88.165 ;
        RECT 93.965 87.995 94.135 88.165 ;
        RECT 94.425 87.995 94.595 88.165 ;
        RECT 94.885 87.995 95.055 88.165 ;
        RECT 95.345 87.995 95.515 88.165 ;
        RECT 95.805 87.995 95.975 88.165 ;
        RECT 96.265 87.995 96.435 88.165 ;
        RECT 96.725 87.995 96.895 88.165 ;
        RECT 97.185 87.995 97.355 88.165 ;
        RECT 97.645 87.995 97.815 88.165 ;
        RECT 98.105 87.995 98.275 88.165 ;
        RECT 98.565 87.995 98.735 88.165 ;
        RECT 99.025 87.995 99.195 88.165 ;
        RECT 99.485 87.995 99.655 88.165 ;
        RECT 99.945 87.995 100.115 88.165 ;
        RECT 100.405 87.995 100.575 88.165 ;
        RECT 100.865 87.995 101.035 88.165 ;
        RECT 101.325 87.995 101.495 88.165 ;
        RECT 101.785 87.995 101.955 88.165 ;
        RECT 102.245 87.995 102.415 88.165 ;
        RECT 102.705 87.995 102.875 88.165 ;
        RECT 103.165 87.995 103.335 88.165 ;
        RECT 103.625 87.995 103.795 88.165 ;
        RECT 104.085 87.995 104.255 88.165 ;
        RECT 104.545 87.995 104.715 88.165 ;
        RECT 105.005 87.995 105.175 88.165 ;
        RECT 105.465 87.995 105.635 88.165 ;
        RECT 105.925 87.995 106.095 88.165 ;
        RECT 106.385 87.995 106.555 88.165 ;
        RECT 106.845 87.995 107.015 88.165 ;
        RECT 107.305 87.995 107.475 88.165 ;
        RECT 107.765 87.995 107.935 88.165 ;
        RECT 108.225 87.995 108.395 88.165 ;
        RECT 108.685 87.995 108.855 88.165 ;
        RECT 109.145 87.995 109.315 88.165 ;
        RECT 109.605 87.995 109.775 88.165 ;
        RECT 110.065 87.995 110.235 88.165 ;
        RECT 110.525 87.995 110.695 88.165 ;
        RECT 110.985 87.995 111.155 88.165 ;
        RECT 111.445 87.995 111.615 88.165 ;
        RECT 111.905 87.995 112.075 88.165 ;
        RECT 112.365 87.995 112.535 88.165 ;
        RECT 112.825 87.995 112.995 88.165 ;
        RECT 113.285 87.995 113.455 88.165 ;
        RECT 113.745 87.995 113.915 88.165 ;
        RECT 114.205 87.995 114.375 88.165 ;
        RECT 114.665 87.995 114.835 88.165 ;
        RECT 115.125 87.995 115.295 88.165 ;
        RECT 115.585 87.995 115.755 88.165 ;
        RECT 116.045 87.995 116.215 88.165 ;
        RECT 116.505 87.995 116.675 88.165 ;
        RECT 116.965 87.995 117.135 88.165 ;
        RECT 117.425 87.995 117.595 88.165 ;
        RECT 117.885 87.995 118.055 88.165 ;
        RECT 118.345 87.995 118.515 88.165 ;
        RECT 118.805 87.995 118.975 88.165 ;
        RECT 119.265 87.995 119.435 88.165 ;
        RECT 119.725 87.995 119.895 88.165 ;
        RECT 120.185 87.995 120.355 88.165 ;
        RECT 120.645 87.995 120.815 88.165 ;
        RECT 121.105 87.995 121.275 88.165 ;
        RECT 121.565 87.995 121.735 88.165 ;
        RECT 122.025 87.995 122.195 88.165 ;
        RECT 122.485 87.995 122.655 88.165 ;
        RECT 122.945 87.995 123.115 88.165 ;
        RECT 123.405 87.995 123.575 88.165 ;
        RECT 123.865 87.995 124.035 88.165 ;
        RECT 124.325 87.995 124.495 88.165 ;
        RECT 124.785 87.995 124.955 88.165 ;
        RECT 125.245 87.995 125.415 88.165 ;
        RECT 125.705 87.995 125.875 88.165 ;
        RECT 126.165 87.995 126.335 88.165 ;
        RECT 126.625 87.995 126.795 88.165 ;
        RECT 127.085 87.995 127.255 88.165 ;
        RECT 127.545 87.995 127.715 88.165 ;
        RECT 128.005 87.995 128.175 88.165 ;
        RECT 128.465 87.995 128.635 88.165 ;
        RECT 128.925 87.995 129.095 88.165 ;
        RECT 129.385 87.995 129.555 88.165 ;
        RECT 129.845 87.995 130.015 88.165 ;
        RECT 130.305 87.995 130.475 88.165 ;
        RECT 130.765 87.995 130.935 88.165 ;
        RECT 131.225 87.995 131.395 88.165 ;
        RECT 131.685 87.995 131.855 88.165 ;
        RECT 132.145 87.995 132.315 88.165 ;
        RECT 132.605 87.995 132.775 88.165 ;
        RECT 133.065 87.995 133.235 88.165 ;
        RECT 133.525 87.995 133.695 88.165 ;
        RECT 133.985 87.995 134.155 88.165 ;
        RECT 45.665 82.555 45.835 82.725 ;
        RECT 46.125 82.555 46.295 82.725 ;
        RECT 46.585 82.555 46.755 82.725 ;
        RECT 47.045 82.555 47.215 82.725 ;
        RECT 47.505 82.555 47.675 82.725 ;
        RECT 47.965 82.555 48.135 82.725 ;
        RECT 48.425 82.555 48.595 82.725 ;
        RECT 48.885 82.555 49.055 82.725 ;
        RECT 49.345 82.555 49.515 82.725 ;
        RECT 49.805 82.555 49.975 82.725 ;
        RECT 50.265 82.555 50.435 82.725 ;
        RECT 50.725 82.555 50.895 82.725 ;
        RECT 51.185 82.555 51.355 82.725 ;
        RECT 51.645 82.555 51.815 82.725 ;
        RECT 52.105 82.555 52.275 82.725 ;
        RECT 52.565 82.555 52.735 82.725 ;
        RECT 53.025 82.555 53.195 82.725 ;
        RECT 53.485 82.555 53.655 82.725 ;
        RECT 53.945 82.555 54.115 82.725 ;
        RECT 54.405 82.555 54.575 82.725 ;
        RECT 54.865 82.555 55.035 82.725 ;
        RECT 55.325 82.555 55.495 82.725 ;
        RECT 55.785 82.555 55.955 82.725 ;
        RECT 56.245 82.555 56.415 82.725 ;
        RECT 56.705 82.555 56.875 82.725 ;
        RECT 57.165 82.555 57.335 82.725 ;
        RECT 57.625 82.555 57.795 82.725 ;
        RECT 58.085 82.555 58.255 82.725 ;
        RECT 58.545 82.555 58.715 82.725 ;
        RECT 59.005 82.555 59.175 82.725 ;
        RECT 59.465 82.555 59.635 82.725 ;
        RECT 59.925 82.555 60.095 82.725 ;
        RECT 60.385 82.555 60.555 82.725 ;
        RECT 60.845 82.555 61.015 82.725 ;
        RECT 61.305 82.555 61.475 82.725 ;
        RECT 61.765 82.555 61.935 82.725 ;
        RECT 62.225 82.555 62.395 82.725 ;
        RECT 62.685 82.555 62.855 82.725 ;
        RECT 63.145 82.555 63.315 82.725 ;
        RECT 63.605 82.555 63.775 82.725 ;
        RECT 64.065 82.555 64.235 82.725 ;
        RECT 64.525 82.555 64.695 82.725 ;
        RECT 64.985 82.555 65.155 82.725 ;
        RECT 65.445 82.555 65.615 82.725 ;
        RECT 65.905 82.555 66.075 82.725 ;
        RECT 66.365 82.555 66.535 82.725 ;
        RECT 66.825 82.555 66.995 82.725 ;
        RECT 67.285 82.555 67.455 82.725 ;
        RECT 67.745 82.555 67.915 82.725 ;
        RECT 68.205 82.555 68.375 82.725 ;
        RECT 68.665 82.555 68.835 82.725 ;
        RECT 69.125 82.555 69.295 82.725 ;
        RECT 69.585 82.555 69.755 82.725 ;
        RECT 70.045 82.555 70.215 82.725 ;
        RECT 70.505 82.555 70.675 82.725 ;
        RECT 70.965 82.555 71.135 82.725 ;
        RECT 71.425 82.555 71.595 82.725 ;
        RECT 71.885 82.555 72.055 82.725 ;
        RECT 72.345 82.555 72.515 82.725 ;
        RECT 72.805 82.555 72.975 82.725 ;
        RECT 73.265 82.555 73.435 82.725 ;
        RECT 73.725 82.555 73.895 82.725 ;
        RECT 74.185 82.555 74.355 82.725 ;
        RECT 74.645 82.555 74.815 82.725 ;
        RECT 75.105 82.555 75.275 82.725 ;
        RECT 75.565 82.555 75.735 82.725 ;
        RECT 76.025 82.555 76.195 82.725 ;
        RECT 76.485 82.555 76.655 82.725 ;
        RECT 76.945 82.555 77.115 82.725 ;
        RECT 77.405 82.555 77.575 82.725 ;
        RECT 77.865 82.555 78.035 82.725 ;
        RECT 78.325 82.555 78.495 82.725 ;
        RECT 78.785 82.555 78.955 82.725 ;
        RECT 79.245 82.555 79.415 82.725 ;
        RECT 79.705 82.555 79.875 82.725 ;
        RECT 80.165 82.555 80.335 82.725 ;
        RECT 80.625 82.555 80.795 82.725 ;
        RECT 81.085 82.555 81.255 82.725 ;
        RECT 81.545 82.555 81.715 82.725 ;
        RECT 82.005 82.555 82.175 82.725 ;
        RECT 82.465 82.555 82.635 82.725 ;
        RECT 82.925 82.555 83.095 82.725 ;
        RECT 83.385 82.555 83.555 82.725 ;
        RECT 83.845 82.555 84.015 82.725 ;
        RECT 84.305 82.555 84.475 82.725 ;
        RECT 84.765 82.555 84.935 82.725 ;
        RECT 85.225 82.555 85.395 82.725 ;
        RECT 85.685 82.555 85.855 82.725 ;
        RECT 86.145 82.555 86.315 82.725 ;
        RECT 86.605 82.555 86.775 82.725 ;
        RECT 87.065 82.555 87.235 82.725 ;
        RECT 87.525 82.555 87.695 82.725 ;
        RECT 87.985 82.555 88.155 82.725 ;
        RECT 88.445 82.555 88.615 82.725 ;
        RECT 88.905 82.555 89.075 82.725 ;
        RECT 89.365 82.555 89.535 82.725 ;
        RECT 89.825 82.555 89.995 82.725 ;
        RECT 90.285 82.555 90.455 82.725 ;
        RECT 90.745 82.555 90.915 82.725 ;
        RECT 91.205 82.555 91.375 82.725 ;
        RECT 91.665 82.555 91.835 82.725 ;
        RECT 92.125 82.555 92.295 82.725 ;
        RECT 92.585 82.555 92.755 82.725 ;
        RECT 93.045 82.555 93.215 82.725 ;
        RECT 93.505 82.555 93.675 82.725 ;
        RECT 93.965 82.555 94.135 82.725 ;
        RECT 94.425 82.555 94.595 82.725 ;
        RECT 94.885 82.555 95.055 82.725 ;
        RECT 95.345 82.555 95.515 82.725 ;
        RECT 95.805 82.555 95.975 82.725 ;
        RECT 96.265 82.555 96.435 82.725 ;
        RECT 96.725 82.555 96.895 82.725 ;
        RECT 97.185 82.555 97.355 82.725 ;
        RECT 97.645 82.555 97.815 82.725 ;
        RECT 98.105 82.555 98.275 82.725 ;
        RECT 98.565 82.555 98.735 82.725 ;
        RECT 99.025 82.555 99.195 82.725 ;
        RECT 99.485 82.555 99.655 82.725 ;
        RECT 99.945 82.555 100.115 82.725 ;
        RECT 100.405 82.555 100.575 82.725 ;
        RECT 100.865 82.555 101.035 82.725 ;
        RECT 101.325 82.555 101.495 82.725 ;
        RECT 101.785 82.555 101.955 82.725 ;
        RECT 102.245 82.555 102.415 82.725 ;
        RECT 102.705 82.555 102.875 82.725 ;
        RECT 103.165 82.555 103.335 82.725 ;
        RECT 103.625 82.555 103.795 82.725 ;
        RECT 104.085 82.555 104.255 82.725 ;
        RECT 104.545 82.555 104.715 82.725 ;
        RECT 105.005 82.555 105.175 82.725 ;
        RECT 105.465 82.555 105.635 82.725 ;
        RECT 105.925 82.555 106.095 82.725 ;
        RECT 106.385 82.555 106.555 82.725 ;
        RECT 106.845 82.555 107.015 82.725 ;
        RECT 107.305 82.555 107.475 82.725 ;
        RECT 107.765 82.555 107.935 82.725 ;
        RECT 108.225 82.555 108.395 82.725 ;
        RECT 108.685 82.555 108.855 82.725 ;
        RECT 109.145 82.555 109.315 82.725 ;
        RECT 109.605 82.555 109.775 82.725 ;
        RECT 110.065 82.555 110.235 82.725 ;
        RECT 110.525 82.555 110.695 82.725 ;
        RECT 110.985 82.555 111.155 82.725 ;
        RECT 111.445 82.555 111.615 82.725 ;
        RECT 111.905 82.555 112.075 82.725 ;
        RECT 112.365 82.555 112.535 82.725 ;
        RECT 112.825 82.555 112.995 82.725 ;
        RECT 113.285 82.555 113.455 82.725 ;
        RECT 113.745 82.555 113.915 82.725 ;
        RECT 114.205 82.555 114.375 82.725 ;
        RECT 114.665 82.555 114.835 82.725 ;
        RECT 115.125 82.555 115.295 82.725 ;
        RECT 115.585 82.555 115.755 82.725 ;
        RECT 116.045 82.555 116.215 82.725 ;
        RECT 116.505 82.555 116.675 82.725 ;
        RECT 116.965 82.555 117.135 82.725 ;
        RECT 117.425 82.555 117.595 82.725 ;
        RECT 117.885 82.555 118.055 82.725 ;
        RECT 118.345 82.555 118.515 82.725 ;
        RECT 118.805 82.555 118.975 82.725 ;
        RECT 119.265 82.555 119.435 82.725 ;
        RECT 119.725 82.555 119.895 82.725 ;
        RECT 120.185 82.555 120.355 82.725 ;
        RECT 120.645 82.555 120.815 82.725 ;
        RECT 121.105 82.555 121.275 82.725 ;
        RECT 121.565 82.555 121.735 82.725 ;
        RECT 122.025 82.555 122.195 82.725 ;
        RECT 122.485 82.555 122.655 82.725 ;
        RECT 122.945 82.555 123.115 82.725 ;
        RECT 123.405 82.555 123.575 82.725 ;
        RECT 123.865 82.555 124.035 82.725 ;
        RECT 124.325 82.555 124.495 82.725 ;
        RECT 124.785 82.555 124.955 82.725 ;
        RECT 125.245 82.555 125.415 82.725 ;
        RECT 125.705 82.555 125.875 82.725 ;
        RECT 126.165 82.555 126.335 82.725 ;
        RECT 126.625 82.555 126.795 82.725 ;
        RECT 127.085 82.555 127.255 82.725 ;
        RECT 127.545 82.555 127.715 82.725 ;
        RECT 128.005 82.555 128.175 82.725 ;
        RECT 128.465 82.555 128.635 82.725 ;
        RECT 128.925 82.555 129.095 82.725 ;
        RECT 129.385 82.555 129.555 82.725 ;
        RECT 129.845 82.555 130.015 82.725 ;
        RECT 130.305 82.555 130.475 82.725 ;
        RECT 130.765 82.555 130.935 82.725 ;
        RECT 131.225 82.555 131.395 82.725 ;
        RECT 131.685 82.555 131.855 82.725 ;
        RECT 132.145 82.555 132.315 82.725 ;
        RECT 132.605 82.555 132.775 82.725 ;
        RECT 133.065 82.555 133.235 82.725 ;
        RECT 133.525 82.555 133.695 82.725 ;
        RECT 133.985 82.555 134.155 82.725 ;
        RECT 45.665 77.115 45.835 77.285 ;
        RECT 46.125 77.115 46.295 77.285 ;
        RECT 46.585 77.115 46.755 77.285 ;
        RECT 47.045 77.115 47.215 77.285 ;
        RECT 47.505 77.115 47.675 77.285 ;
        RECT 47.965 77.115 48.135 77.285 ;
        RECT 48.425 77.115 48.595 77.285 ;
        RECT 48.885 77.115 49.055 77.285 ;
        RECT 49.345 77.115 49.515 77.285 ;
        RECT 49.805 77.115 49.975 77.285 ;
        RECT 50.265 77.115 50.435 77.285 ;
        RECT 50.725 77.115 50.895 77.285 ;
        RECT 51.185 77.115 51.355 77.285 ;
        RECT 51.645 77.115 51.815 77.285 ;
        RECT 52.105 77.115 52.275 77.285 ;
        RECT 52.565 77.115 52.735 77.285 ;
        RECT 53.025 77.115 53.195 77.285 ;
        RECT 53.485 77.115 53.655 77.285 ;
        RECT 53.945 77.115 54.115 77.285 ;
        RECT 54.405 77.115 54.575 77.285 ;
        RECT 54.865 77.115 55.035 77.285 ;
        RECT 55.325 77.115 55.495 77.285 ;
        RECT 55.785 77.115 55.955 77.285 ;
        RECT 56.245 77.115 56.415 77.285 ;
        RECT 56.705 77.115 56.875 77.285 ;
        RECT 57.165 77.115 57.335 77.285 ;
        RECT 57.625 77.115 57.795 77.285 ;
        RECT 58.085 77.115 58.255 77.285 ;
        RECT 58.545 77.115 58.715 77.285 ;
        RECT 59.005 77.115 59.175 77.285 ;
        RECT 59.465 77.115 59.635 77.285 ;
        RECT 59.925 77.115 60.095 77.285 ;
        RECT 60.385 77.115 60.555 77.285 ;
        RECT 60.845 77.115 61.015 77.285 ;
        RECT 61.305 77.115 61.475 77.285 ;
        RECT 61.765 77.115 61.935 77.285 ;
        RECT 62.225 77.115 62.395 77.285 ;
        RECT 62.685 77.115 62.855 77.285 ;
        RECT 63.145 77.115 63.315 77.285 ;
        RECT 63.605 77.115 63.775 77.285 ;
        RECT 64.065 77.115 64.235 77.285 ;
        RECT 64.525 77.115 64.695 77.285 ;
        RECT 64.985 77.115 65.155 77.285 ;
        RECT 65.445 77.115 65.615 77.285 ;
        RECT 65.905 77.115 66.075 77.285 ;
        RECT 66.365 77.115 66.535 77.285 ;
        RECT 66.825 77.115 66.995 77.285 ;
        RECT 67.285 77.115 67.455 77.285 ;
        RECT 67.745 77.115 67.915 77.285 ;
        RECT 68.205 77.115 68.375 77.285 ;
        RECT 68.665 77.115 68.835 77.285 ;
        RECT 69.125 77.115 69.295 77.285 ;
        RECT 69.585 77.115 69.755 77.285 ;
        RECT 70.045 77.115 70.215 77.285 ;
        RECT 70.505 77.115 70.675 77.285 ;
        RECT 70.965 77.115 71.135 77.285 ;
        RECT 71.425 77.115 71.595 77.285 ;
        RECT 71.885 77.115 72.055 77.285 ;
        RECT 72.345 77.115 72.515 77.285 ;
        RECT 72.805 77.115 72.975 77.285 ;
        RECT 73.265 77.115 73.435 77.285 ;
        RECT 73.725 77.115 73.895 77.285 ;
        RECT 74.185 77.115 74.355 77.285 ;
        RECT 74.645 77.115 74.815 77.285 ;
        RECT 75.105 77.115 75.275 77.285 ;
        RECT 75.565 77.115 75.735 77.285 ;
        RECT 76.025 77.115 76.195 77.285 ;
        RECT 76.485 77.115 76.655 77.285 ;
        RECT 76.945 77.115 77.115 77.285 ;
        RECT 77.405 77.115 77.575 77.285 ;
        RECT 77.865 77.115 78.035 77.285 ;
        RECT 78.325 77.115 78.495 77.285 ;
        RECT 78.785 77.115 78.955 77.285 ;
        RECT 79.245 77.115 79.415 77.285 ;
        RECT 79.705 77.115 79.875 77.285 ;
        RECT 80.165 77.115 80.335 77.285 ;
        RECT 80.625 77.115 80.795 77.285 ;
        RECT 81.085 77.115 81.255 77.285 ;
        RECT 81.545 77.115 81.715 77.285 ;
        RECT 82.005 77.115 82.175 77.285 ;
        RECT 82.465 77.115 82.635 77.285 ;
        RECT 82.925 77.115 83.095 77.285 ;
        RECT 83.385 77.115 83.555 77.285 ;
        RECT 83.845 77.115 84.015 77.285 ;
        RECT 84.305 77.115 84.475 77.285 ;
        RECT 84.765 77.115 84.935 77.285 ;
        RECT 85.225 77.115 85.395 77.285 ;
        RECT 85.685 77.115 85.855 77.285 ;
        RECT 86.145 77.115 86.315 77.285 ;
        RECT 86.605 77.115 86.775 77.285 ;
        RECT 87.065 77.115 87.235 77.285 ;
        RECT 87.525 77.115 87.695 77.285 ;
        RECT 87.985 77.115 88.155 77.285 ;
        RECT 88.445 77.115 88.615 77.285 ;
        RECT 88.905 77.115 89.075 77.285 ;
        RECT 89.365 77.115 89.535 77.285 ;
        RECT 89.825 77.115 89.995 77.285 ;
        RECT 90.285 77.115 90.455 77.285 ;
        RECT 90.745 77.115 90.915 77.285 ;
        RECT 91.205 77.115 91.375 77.285 ;
        RECT 91.665 77.115 91.835 77.285 ;
        RECT 92.125 77.115 92.295 77.285 ;
        RECT 92.585 77.115 92.755 77.285 ;
        RECT 93.045 77.115 93.215 77.285 ;
        RECT 93.505 77.115 93.675 77.285 ;
        RECT 93.965 77.115 94.135 77.285 ;
        RECT 94.425 77.115 94.595 77.285 ;
        RECT 94.885 77.115 95.055 77.285 ;
        RECT 95.345 77.115 95.515 77.285 ;
        RECT 95.805 77.115 95.975 77.285 ;
        RECT 96.265 77.115 96.435 77.285 ;
        RECT 96.725 77.115 96.895 77.285 ;
        RECT 97.185 77.115 97.355 77.285 ;
        RECT 97.645 77.115 97.815 77.285 ;
        RECT 98.105 77.115 98.275 77.285 ;
        RECT 98.565 77.115 98.735 77.285 ;
        RECT 99.025 77.115 99.195 77.285 ;
        RECT 99.485 77.115 99.655 77.285 ;
        RECT 99.945 77.115 100.115 77.285 ;
        RECT 100.405 77.115 100.575 77.285 ;
        RECT 100.865 77.115 101.035 77.285 ;
        RECT 101.325 77.115 101.495 77.285 ;
        RECT 101.785 77.115 101.955 77.285 ;
        RECT 102.245 77.115 102.415 77.285 ;
        RECT 102.705 77.115 102.875 77.285 ;
        RECT 103.165 77.115 103.335 77.285 ;
        RECT 103.625 77.115 103.795 77.285 ;
        RECT 104.085 77.115 104.255 77.285 ;
        RECT 104.545 77.115 104.715 77.285 ;
        RECT 105.005 77.115 105.175 77.285 ;
        RECT 105.465 77.115 105.635 77.285 ;
        RECT 105.925 77.115 106.095 77.285 ;
        RECT 106.385 77.115 106.555 77.285 ;
        RECT 106.845 77.115 107.015 77.285 ;
        RECT 107.305 77.115 107.475 77.285 ;
        RECT 107.765 77.115 107.935 77.285 ;
        RECT 108.225 77.115 108.395 77.285 ;
        RECT 108.685 77.115 108.855 77.285 ;
        RECT 109.145 77.115 109.315 77.285 ;
        RECT 109.605 77.115 109.775 77.285 ;
        RECT 110.065 77.115 110.235 77.285 ;
        RECT 110.525 77.115 110.695 77.285 ;
        RECT 110.985 77.115 111.155 77.285 ;
        RECT 111.445 77.115 111.615 77.285 ;
        RECT 111.905 77.115 112.075 77.285 ;
        RECT 112.365 77.115 112.535 77.285 ;
        RECT 112.825 77.115 112.995 77.285 ;
        RECT 113.285 77.115 113.455 77.285 ;
        RECT 113.745 77.115 113.915 77.285 ;
        RECT 114.205 77.115 114.375 77.285 ;
        RECT 114.665 77.115 114.835 77.285 ;
        RECT 115.125 77.115 115.295 77.285 ;
        RECT 115.585 77.115 115.755 77.285 ;
        RECT 116.045 77.115 116.215 77.285 ;
        RECT 116.505 77.115 116.675 77.285 ;
        RECT 116.965 77.115 117.135 77.285 ;
        RECT 117.425 77.115 117.595 77.285 ;
        RECT 117.885 77.115 118.055 77.285 ;
        RECT 118.345 77.115 118.515 77.285 ;
        RECT 118.805 77.115 118.975 77.285 ;
        RECT 119.265 77.115 119.435 77.285 ;
        RECT 119.725 77.115 119.895 77.285 ;
        RECT 120.185 77.115 120.355 77.285 ;
        RECT 120.645 77.115 120.815 77.285 ;
        RECT 121.105 77.115 121.275 77.285 ;
        RECT 121.565 77.115 121.735 77.285 ;
        RECT 122.025 77.115 122.195 77.285 ;
        RECT 122.485 77.115 122.655 77.285 ;
        RECT 122.945 77.115 123.115 77.285 ;
        RECT 123.405 77.115 123.575 77.285 ;
        RECT 123.865 77.115 124.035 77.285 ;
        RECT 124.325 77.115 124.495 77.285 ;
        RECT 124.785 77.115 124.955 77.285 ;
        RECT 125.245 77.115 125.415 77.285 ;
        RECT 125.705 77.115 125.875 77.285 ;
        RECT 126.165 77.115 126.335 77.285 ;
        RECT 126.625 77.115 126.795 77.285 ;
        RECT 127.085 77.115 127.255 77.285 ;
        RECT 127.545 77.115 127.715 77.285 ;
        RECT 128.005 77.115 128.175 77.285 ;
        RECT 128.465 77.115 128.635 77.285 ;
        RECT 128.925 77.115 129.095 77.285 ;
        RECT 129.385 77.115 129.555 77.285 ;
        RECT 129.845 77.115 130.015 77.285 ;
        RECT 130.305 77.115 130.475 77.285 ;
        RECT 130.765 77.115 130.935 77.285 ;
        RECT 131.225 77.115 131.395 77.285 ;
        RECT 131.685 77.115 131.855 77.285 ;
        RECT 132.145 77.115 132.315 77.285 ;
        RECT 132.605 77.115 132.775 77.285 ;
        RECT 133.065 77.115 133.235 77.285 ;
        RECT 133.525 77.115 133.695 77.285 ;
        RECT 133.985 77.115 134.155 77.285 ;
        RECT 45.665 71.675 45.835 71.845 ;
        RECT 46.125 71.675 46.295 71.845 ;
        RECT 46.585 71.675 46.755 71.845 ;
        RECT 47.045 71.675 47.215 71.845 ;
        RECT 47.505 71.675 47.675 71.845 ;
        RECT 47.965 71.675 48.135 71.845 ;
        RECT 48.425 71.675 48.595 71.845 ;
        RECT 48.885 71.675 49.055 71.845 ;
        RECT 49.345 71.675 49.515 71.845 ;
        RECT 49.805 71.675 49.975 71.845 ;
        RECT 50.265 71.675 50.435 71.845 ;
        RECT 50.725 71.675 50.895 71.845 ;
        RECT 51.185 71.675 51.355 71.845 ;
        RECT 51.645 71.675 51.815 71.845 ;
        RECT 52.105 71.675 52.275 71.845 ;
        RECT 52.565 71.675 52.735 71.845 ;
        RECT 53.025 71.675 53.195 71.845 ;
        RECT 53.485 71.675 53.655 71.845 ;
        RECT 53.945 71.675 54.115 71.845 ;
        RECT 54.405 71.675 54.575 71.845 ;
        RECT 54.865 71.675 55.035 71.845 ;
        RECT 55.325 71.675 55.495 71.845 ;
        RECT 55.785 71.675 55.955 71.845 ;
        RECT 56.245 71.675 56.415 71.845 ;
        RECT 56.705 71.675 56.875 71.845 ;
        RECT 57.165 71.675 57.335 71.845 ;
        RECT 57.625 71.675 57.795 71.845 ;
        RECT 58.085 71.675 58.255 71.845 ;
        RECT 58.545 71.675 58.715 71.845 ;
        RECT 59.005 71.675 59.175 71.845 ;
        RECT 59.465 71.675 59.635 71.845 ;
        RECT 59.925 71.675 60.095 71.845 ;
        RECT 60.385 71.675 60.555 71.845 ;
        RECT 60.845 71.675 61.015 71.845 ;
        RECT 61.305 71.675 61.475 71.845 ;
        RECT 61.765 71.675 61.935 71.845 ;
        RECT 62.225 71.675 62.395 71.845 ;
        RECT 62.685 71.675 62.855 71.845 ;
        RECT 63.145 71.675 63.315 71.845 ;
        RECT 63.605 71.675 63.775 71.845 ;
        RECT 64.065 71.675 64.235 71.845 ;
        RECT 64.525 71.675 64.695 71.845 ;
        RECT 64.985 71.675 65.155 71.845 ;
        RECT 65.445 71.675 65.615 71.845 ;
        RECT 65.905 71.675 66.075 71.845 ;
        RECT 66.365 71.675 66.535 71.845 ;
        RECT 66.825 71.675 66.995 71.845 ;
        RECT 67.285 71.675 67.455 71.845 ;
        RECT 67.745 71.675 67.915 71.845 ;
        RECT 68.205 71.675 68.375 71.845 ;
        RECT 68.665 71.675 68.835 71.845 ;
        RECT 69.125 71.675 69.295 71.845 ;
        RECT 69.585 71.675 69.755 71.845 ;
        RECT 70.045 71.675 70.215 71.845 ;
        RECT 70.505 71.675 70.675 71.845 ;
        RECT 70.965 71.675 71.135 71.845 ;
        RECT 71.425 71.675 71.595 71.845 ;
        RECT 71.885 71.675 72.055 71.845 ;
        RECT 72.345 71.675 72.515 71.845 ;
        RECT 72.805 71.675 72.975 71.845 ;
        RECT 73.265 71.675 73.435 71.845 ;
        RECT 73.725 71.675 73.895 71.845 ;
        RECT 74.185 71.675 74.355 71.845 ;
        RECT 74.645 71.675 74.815 71.845 ;
        RECT 75.105 71.675 75.275 71.845 ;
        RECT 75.565 71.675 75.735 71.845 ;
        RECT 76.025 71.675 76.195 71.845 ;
        RECT 76.485 71.675 76.655 71.845 ;
        RECT 76.945 71.675 77.115 71.845 ;
        RECT 77.405 71.675 77.575 71.845 ;
        RECT 77.865 71.675 78.035 71.845 ;
        RECT 78.325 71.675 78.495 71.845 ;
        RECT 78.785 71.675 78.955 71.845 ;
        RECT 79.245 71.675 79.415 71.845 ;
        RECT 79.705 71.675 79.875 71.845 ;
        RECT 80.165 71.675 80.335 71.845 ;
        RECT 80.625 71.675 80.795 71.845 ;
        RECT 81.085 71.675 81.255 71.845 ;
        RECT 81.545 71.675 81.715 71.845 ;
        RECT 82.005 71.675 82.175 71.845 ;
        RECT 82.465 71.675 82.635 71.845 ;
        RECT 82.925 71.675 83.095 71.845 ;
        RECT 83.385 71.675 83.555 71.845 ;
        RECT 83.845 71.675 84.015 71.845 ;
        RECT 84.305 71.675 84.475 71.845 ;
        RECT 84.765 71.675 84.935 71.845 ;
        RECT 85.225 71.675 85.395 71.845 ;
        RECT 85.685 71.675 85.855 71.845 ;
        RECT 86.145 71.675 86.315 71.845 ;
        RECT 86.605 71.675 86.775 71.845 ;
        RECT 87.065 71.675 87.235 71.845 ;
        RECT 87.525 71.675 87.695 71.845 ;
        RECT 87.985 71.675 88.155 71.845 ;
        RECT 88.445 71.675 88.615 71.845 ;
        RECT 88.905 71.675 89.075 71.845 ;
        RECT 89.365 71.675 89.535 71.845 ;
        RECT 89.825 71.675 89.995 71.845 ;
        RECT 90.285 71.675 90.455 71.845 ;
        RECT 90.745 71.675 90.915 71.845 ;
        RECT 91.205 71.675 91.375 71.845 ;
        RECT 91.665 71.675 91.835 71.845 ;
        RECT 92.125 71.675 92.295 71.845 ;
        RECT 92.585 71.675 92.755 71.845 ;
        RECT 93.045 71.675 93.215 71.845 ;
        RECT 93.505 71.675 93.675 71.845 ;
        RECT 93.965 71.675 94.135 71.845 ;
        RECT 94.425 71.675 94.595 71.845 ;
        RECT 94.885 71.675 95.055 71.845 ;
        RECT 95.345 71.675 95.515 71.845 ;
        RECT 95.805 71.675 95.975 71.845 ;
        RECT 96.265 71.675 96.435 71.845 ;
        RECT 96.725 71.675 96.895 71.845 ;
        RECT 97.185 71.675 97.355 71.845 ;
        RECT 97.645 71.675 97.815 71.845 ;
        RECT 98.105 71.675 98.275 71.845 ;
        RECT 98.565 71.675 98.735 71.845 ;
        RECT 99.025 71.675 99.195 71.845 ;
        RECT 99.485 71.675 99.655 71.845 ;
        RECT 99.945 71.675 100.115 71.845 ;
        RECT 100.405 71.675 100.575 71.845 ;
        RECT 100.865 71.675 101.035 71.845 ;
        RECT 101.325 71.675 101.495 71.845 ;
        RECT 101.785 71.675 101.955 71.845 ;
        RECT 102.245 71.675 102.415 71.845 ;
        RECT 102.705 71.675 102.875 71.845 ;
        RECT 103.165 71.675 103.335 71.845 ;
        RECT 103.625 71.675 103.795 71.845 ;
        RECT 104.085 71.675 104.255 71.845 ;
        RECT 104.545 71.675 104.715 71.845 ;
        RECT 105.005 71.675 105.175 71.845 ;
        RECT 105.465 71.675 105.635 71.845 ;
        RECT 105.925 71.675 106.095 71.845 ;
        RECT 106.385 71.675 106.555 71.845 ;
        RECT 106.845 71.675 107.015 71.845 ;
        RECT 107.305 71.675 107.475 71.845 ;
        RECT 107.765 71.675 107.935 71.845 ;
        RECT 108.225 71.675 108.395 71.845 ;
        RECT 108.685 71.675 108.855 71.845 ;
        RECT 109.145 71.675 109.315 71.845 ;
        RECT 109.605 71.675 109.775 71.845 ;
        RECT 110.065 71.675 110.235 71.845 ;
        RECT 110.525 71.675 110.695 71.845 ;
        RECT 110.985 71.675 111.155 71.845 ;
        RECT 111.445 71.675 111.615 71.845 ;
        RECT 111.905 71.675 112.075 71.845 ;
        RECT 112.365 71.675 112.535 71.845 ;
        RECT 112.825 71.675 112.995 71.845 ;
        RECT 113.285 71.675 113.455 71.845 ;
        RECT 113.745 71.675 113.915 71.845 ;
        RECT 114.205 71.675 114.375 71.845 ;
        RECT 114.665 71.675 114.835 71.845 ;
        RECT 115.125 71.675 115.295 71.845 ;
        RECT 115.585 71.675 115.755 71.845 ;
        RECT 116.045 71.675 116.215 71.845 ;
        RECT 116.505 71.675 116.675 71.845 ;
        RECT 116.965 71.675 117.135 71.845 ;
        RECT 117.425 71.675 117.595 71.845 ;
        RECT 117.885 71.675 118.055 71.845 ;
        RECT 118.345 71.675 118.515 71.845 ;
        RECT 118.805 71.675 118.975 71.845 ;
        RECT 119.265 71.675 119.435 71.845 ;
        RECT 119.725 71.675 119.895 71.845 ;
        RECT 120.185 71.675 120.355 71.845 ;
        RECT 120.645 71.675 120.815 71.845 ;
        RECT 121.105 71.675 121.275 71.845 ;
        RECT 121.565 71.675 121.735 71.845 ;
        RECT 122.025 71.675 122.195 71.845 ;
        RECT 122.485 71.675 122.655 71.845 ;
        RECT 122.945 71.675 123.115 71.845 ;
        RECT 123.405 71.675 123.575 71.845 ;
        RECT 123.865 71.675 124.035 71.845 ;
        RECT 124.325 71.675 124.495 71.845 ;
        RECT 124.785 71.675 124.955 71.845 ;
        RECT 125.245 71.675 125.415 71.845 ;
        RECT 125.705 71.675 125.875 71.845 ;
        RECT 126.165 71.675 126.335 71.845 ;
        RECT 126.625 71.675 126.795 71.845 ;
        RECT 127.085 71.675 127.255 71.845 ;
        RECT 127.545 71.675 127.715 71.845 ;
        RECT 128.005 71.675 128.175 71.845 ;
        RECT 128.465 71.675 128.635 71.845 ;
        RECT 128.925 71.675 129.095 71.845 ;
        RECT 129.385 71.675 129.555 71.845 ;
        RECT 129.845 71.675 130.015 71.845 ;
        RECT 130.305 71.675 130.475 71.845 ;
        RECT 130.765 71.675 130.935 71.845 ;
        RECT 131.225 71.675 131.395 71.845 ;
        RECT 131.685 71.675 131.855 71.845 ;
        RECT 132.145 71.675 132.315 71.845 ;
        RECT 132.605 71.675 132.775 71.845 ;
        RECT 133.065 71.675 133.235 71.845 ;
        RECT 133.525 71.675 133.695 71.845 ;
        RECT 133.985 71.675 134.155 71.845 ;
        RECT 45.665 66.235 45.835 66.405 ;
        RECT 46.125 66.235 46.295 66.405 ;
        RECT 46.585 66.235 46.755 66.405 ;
        RECT 47.045 66.235 47.215 66.405 ;
        RECT 47.505 66.235 47.675 66.405 ;
        RECT 47.965 66.235 48.135 66.405 ;
        RECT 48.425 66.235 48.595 66.405 ;
        RECT 48.885 66.235 49.055 66.405 ;
        RECT 49.345 66.235 49.515 66.405 ;
        RECT 49.805 66.235 49.975 66.405 ;
        RECT 50.265 66.235 50.435 66.405 ;
        RECT 50.725 66.235 50.895 66.405 ;
        RECT 51.185 66.235 51.355 66.405 ;
        RECT 51.645 66.235 51.815 66.405 ;
        RECT 52.105 66.235 52.275 66.405 ;
        RECT 52.565 66.235 52.735 66.405 ;
        RECT 53.025 66.235 53.195 66.405 ;
        RECT 53.485 66.235 53.655 66.405 ;
        RECT 53.945 66.235 54.115 66.405 ;
        RECT 54.405 66.235 54.575 66.405 ;
        RECT 54.865 66.235 55.035 66.405 ;
        RECT 55.325 66.235 55.495 66.405 ;
        RECT 55.785 66.235 55.955 66.405 ;
        RECT 56.245 66.235 56.415 66.405 ;
        RECT 56.705 66.235 56.875 66.405 ;
        RECT 57.165 66.235 57.335 66.405 ;
        RECT 57.625 66.235 57.795 66.405 ;
        RECT 58.085 66.235 58.255 66.405 ;
        RECT 58.545 66.235 58.715 66.405 ;
        RECT 59.005 66.235 59.175 66.405 ;
        RECT 59.465 66.235 59.635 66.405 ;
        RECT 59.925 66.235 60.095 66.405 ;
        RECT 60.385 66.235 60.555 66.405 ;
        RECT 60.845 66.235 61.015 66.405 ;
        RECT 61.305 66.235 61.475 66.405 ;
        RECT 61.765 66.235 61.935 66.405 ;
        RECT 62.225 66.235 62.395 66.405 ;
        RECT 62.685 66.235 62.855 66.405 ;
        RECT 63.145 66.235 63.315 66.405 ;
        RECT 63.605 66.235 63.775 66.405 ;
        RECT 64.065 66.235 64.235 66.405 ;
        RECT 64.525 66.235 64.695 66.405 ;
        RECT 64.985 66.235 65.155 66.405 ;
        RECT 65.445 66.235 65.615 66.405 ;
        RECT 65.905 66.235 66.075 66.405 ;
        RECT 66.365 66.235 66.535 66.405 ;
        RECT 66.825 66.235 66.995 66.405 ;
        RECT 67.285 66.235 67.455 66.405 ;
        RECT 67.745 66.235 67.915 66.405 ;
        RECT 68.205 66.235 68.375 66.405 ;
        RECT 68.665 66.235 68.835 66.405 ;
        RECT 69.125 66.235 69.295 66.405 ;
        RECT 69.585 66.235 69.755 66.405 ;
        RECT 70.045 66.235 70.215 66.405 ;
        RECT 70.505 66.235 70.675 66.405 ;
        RECT 70.965 66.235 71.135 66.405 ;
        RECT 71.425 66.235 71.595 66.405 ;
        RECT 71.885 66.235 72.055 66.405 ;
        RECT 72.345 66.235 72.515 66.405 ;
        RECT 72.805 66.235 72.975 66.405 ;
        RECT 73.265 66.235 73.435 66.405 ;
        RECT 73.725 66.235 73.895 66.405 ;
        RECT 74.185 66.235 74.355 66.405 ;
        RECT 74.645 66.235 74.815 66.405 ;
        RECT 75.105 66.235 75.275 66.405 ;
        RECT 75.565 66.235 75.735 66.405 ;
        RECT 76.025 66.235 76.195 66.405 ;
        RECT 76.485 66.235 76.655 66.405 ;
        RECT 76.945 66.235 77.115 66.405 ;
        RECT 77.405 66.235 77.575 66.405 ;
        RECT 77.865 66.235 78.035 66.405 ;
        RECT 78.325 66.235 78.495 66.405 ;
        RECT 78.785 66.235 78.955 66.405 ;
        RECT 79.245 66.235 79.415 66.405 ;
        RECT 79.705 66.235 79.875 66.405 ;
        RECT 80.165 66.235 80.335 66.405 ;
        RECT 80.625 66.235 80.795 66.405 ;
        RECT 81.085 66.235 81.255 66.405 ;
        RECT 81.545 66.235 81.715 66.405 ;
        RECT 82.005 66.235 82.175 66.405 ;
        RECT 82.465 66.235 82.635 66.405 ;
        RECT 82.925 66.235 83.095 66.405 ;
        RECT 83.385 66.235 83.555 66.405 ;
        RECT 83.845 66.235 84.015 66.405 ;
        RECT 84.305 66.235 84.475 66.405 ;
        RECT 84.765 66.235 84.935 66.405 ;
        RECT 85.225 66.235 85.395 66.405 ;
        RECT 85.685 66.235 85.855 66.405 ;
        RECT 86.145 66.235 86.315 66.405 ;
        RECT 86.605 66.235 86.775 66.405 ;
        RECT 87.065 66.235 87.235 66.405 ;
        RECT 87.525 66.235 87.695 66.405 ;
        RECT 87.985 66.235 88.155 66.405 ;
        RECT 88.445 66.235 88.615 66.405 ;
        RECT 88.905 66.235 89.075 66.405 ;
        RECT 89.365 66.235 89.535 66.405 ;
        RECT 89.825 66.235 89.995 66.405 ;
        RECT 90.285 66.235 90.455 66.405 ;
        RECT 90.745 66.235 90.915 66.405 ;
        RECT 91.205 66.235 91.375 66.405 ;
        RECT 91.665 66.235 91.835 66.405 ;
        RECT 92.125 66.235 92.295 66.405 ;
        RECT 92.585 66.235 92.755 66.405 ;
        RECT 93.045 66.235 93.215 66.405 ;
        RECT 93.505 66.235 93.675 66.405 ;
        RECT 93.965 66.235 94.135 66.405 ;
        RECT 94.425 66.235 94.595 66.405 ;
        RECT 94.885 66.235 95.055 66.405 ;
        RECT 95.345 66.235 95.515 66.405 ;
        RECT 95.805 66.235 95.975 66.405 ;
        RECT 96.265 66.235 96.435 66.405 ;
        RECT 96.725 66.235 96.895 66.405 ;
        RECT 97.185 66.235 97.355 66.405 ;
        RECT 97.645 66.235 97.815 66.405 ;
        RECT 98.105 66.235 98.275 66.405 ;
        RECT 98.565 66.235 98.735 66.405 ;
        RECT 99.025 66.235 99.195 66.405 ;
        RECT 99.485 66.235 99.655 66.405 ;
        RECT 99.945 66.235 100.115 66.405 ;
        RECT 100.405 66.235 100.575 66.405 ;
        RECT 100.865 66.235 101.035 66.405 ;
        RECT 101.325 66.235 101.495 66.405 ;
        RECT 101.785 66.235 101.955 66.405 ;
        RECT 102.245 66.235 102.415 66.405 ;
        RECT 102.705 66.235 102.875 66.405 ;
        RECT 103.165 66.235 103.335 66.405 ;
        RECT 103.625 66.235 103.795 66.405 ;
        RECT 104.085 66.235 104.255 66.405 ;
        RECT 104.545 66.235 104.715 66.405 ;
        RECT 105.005 66.235 105.175 66.405 ;
        RECT 105.465 66.235 105.635 66.405 ;
        RECT 105.925 66.235 106.095 66.405 ;
        RECT 106.385 66.235 106.555 66.405 ;
        RECT 106.845 66.235 107.015 66.405 ;
        RECT 107.305 66.235 107.475 66.405 ;
        RECT 107.765 66.235 107.935 66.405 ;
        RECT 108.225 66.235 108.395 66.405 ;
        RECT 108.685 66.235 108.855 66.405 ;
        RECT 109.145 66.235 109.315 66.405 ;
        RECT 109.605 66.235 109.775 66.405 ;
        RECT 110.065 66.235 110.235 66.405 ;
        RECT 110.525 66.235 110.695 66.405 ;
        RECT 110.985 66.235 111.155 66.405 ;
        RECT 111.445 66.235 111.615 66.405 ;
        RECT 111.905 66.235 112.075 66.405 ;
        RECT 112.365 66.235 112.535 66.405 ;
        RECT 112.825 66.235 112.995 66.405 ;
        RECT 113.285 66.235 113.455 66.405 ;
        RECT 113.745 66.235 113.915 66.405 ;
        RECT 114.205 66.235 114.375 66.405 ;
        RECT 114.665 66.235 114.835 66.405 ;
        RECT 115.125 66.235 115.295 66.405 ;
        RECT 115.585 66.235 115.755 66.405 ;
        RECT 116.045 66.235 116.215 66.405 ;
        RECT 116.505 66.235 116.675 66.405 ;
        RECT 116.965 66.235 117.135 66.405 ;
        RECT 117.425 66.235 117.595 66.405 ;
        RECT 117.885 66.235 118.055 66.405 ;
        RECT 118.345 66.235 118.515 66.405 ;
        RECT 118.805 66.235 118.975 66.405 ;
        RECT 119.265 66.235 119.435 66.405 ;
        RECT 119.725 66.235 119.895 66.405 ;
        RECT 120.185 66.235 120.355 66.405 ;
        RECT 120.645 66.235 120.815 66.405 ;
        RECT 121.105 66.235 121.275 66.405 ;
        RECT 121.565 66.235 121.735 66.405 ;
        RECT 122.025 66.235 122.195 66.405 ;
        RECT 122.485 66.235 122.655 66.405 ;
        RECT 122.945 66.235 123.115 66.405 ;
        RECT 123.405 66.235 123.575 66.405 ;
        RECT 123.865 66.235 124.035 66.405 ;
        RECT 124.325 66.235 124.495 66.405 ;
        RECT 124.785 66.235 124.955 66.405 ;
        RECT 125.245 66.235 125.415 66.405 ;
        RECT 125.705 66.235 125.875 66.405 ;
        RECT 126.165 66.235 126.335 66.405 ;
        RECT 126.625 66.235 126.795 66.405 ;
        RECT 127.085 66.235 127.255 66.405 ;
        RECT 127.545 66.235 127.715 66.405 ;
        RECT 128.005 66.235 128.175 66.405 ;
        RECT 128.465 66.235 128.635 66.405 ;
        RECT 128.925 66.235 129.095 66.405 ;
        RECT 129.385 66.235 129.555 66.405 ;
        RECT 129.845 66.235 130.015 66.405 ;
        RECT 130.305 66.235 130.475 66.405 ;
        RECT 130.765 66.235 130.935 66.405 ;
        RECT 131.225 66.235 131.395 66.405 ;
        RECT 131.685 66.235 131.855 66.405 ;
        RECT 132.145 66.235 132.315 66.405 ;
        RECT 132.605 66.235 132.775 66.405 ;
        RECT 133.065 66.235 133.235 66.405 ;
        RECT 133.525 66.235 133.695 66.405 ;
        RECT 133.985 66.235 134.155 66.405 ;
        RECT 45.665 60.795 45.835 60.965 ;
        RECT 46.125 60.795 46.295 60.965 ;
        RECT 46.585 60.795 46.755 60.965 ;
        RECT 47.045 60.795 47.215 60.965 ;
        RECT 47.505 60.795 47.675 60.965 ;
        RECT 47.965 60.795 48.135 60.965 ;
        RECT 48.425 60.795 48.595 60.965 ;
        RECT 48.885 60.795 49.055 60.965 ;
        RECT 49.345 60.795 49.515 60.965 ;
        RECT 49.805 60.795 49.975 60.965 ;
        RECT 50.265 60.795 50.435 60.965 ;
        RECT 50.725 60.795 50.895 60.965 ;
        RECT 51.185 60.795 51.355 60.965 ;
        RECT 51.645 60.795 51.815 60.965 ;
        RECT 52.105 60.795 52.275 60.965 ;
        RECT 52.565 60.795 52.735 60.965 ;
        RECT 53.025 60.795 53.195 60.965 ;
        RECT 53.485 60.795 53.655 60.965 ;
        RECT 53.945 60.795 54.115 60.965 ;
        RECT 54.405 60.795 54.575 60.965 ;
        RECT 54.865 60.795 55.035 60.965 ;
        RECT 55.325 60.795 55.495 60.965 ;
        RECT 55.785 60.795 55.955 60.965 ;
        RECT 56.245 60.795 56.415 60.965 ;
        RECT 56.705 60.795 56.875 60.965 ;
        RECT 57.165 60.795 57.335 60.965 ;
        RECT 57.625 60.795 57.795 60.965 ;
        RECT 58.085 60.795 58.255 60.965 ;
        RECT 58.545 60.795 58.715 60.965 ;
        RECT 59.005 60.795 59.175 60.965 ;
        RECT 59.465 60.795 59.635 60.965 ;
        RECT 59.925 60.795 60.095 60.965 ;
        RECT 60.385 60.795 60.555 60.965 ;
        RECT 60.845 60.795 61.015 60.965 ;
        RECT 61.305 60.795 61.475 60.965 ;
        RECT 61.765 60.795 61.935 60.965 ;
        RECT 62.225 60.795 62.395 60.965 ;
        RECT 62.685 60.795 62.855 60.965 ;
        RECT 63.145 60.795 63.315 60.965 ;
        RECT 63.605 60.795 63.775 60.965 ;
        RECT 64.065 60.795 64.235 60.965 ;
        RECT 64.525 60.795 64.695 60.965 ;
        RECT 64.985 60.795 65.155 60.965 ;
        RECT 65.445 60.795 65.615 60.965 ;
        RECT 65.905 60.795 66.075 60.965 ;
        RECT 66.365 60.795 66.535 60.965 ;
        RECT 66.825 60.795 66.995 60.965 ;
        RECT 67.285 60.795 67.455 60.965 ;
        RECT 67.745 60.795 67.915 60.965 ;
        RECT 68.205 60.795 68.375 60.965 ;
        RECT 68.665 60.795 68.835 60.965 ;
        RECT 69.125 60.795 69.295 60.965 ;
        RECT 69.585 60.795 69.755 60.965 ;
        RECT 70.045 60.795 70.215 60.965 ;
        RECT 70.505 60.795 70.675 60.965 ;
        RECT 70.965 60.795 71.135 60.965 ;
        RECT 71.425 60.795 71.595 60.965 ;
        RECT 71.885 60.795 72.055 60.965 ;
        RECT 72.345 60.795 72.515 60.965 ;
        RECT 72.805 60.795 72.975 60.965 ;
        RECT 73.265 60.795 73.435 60.965 ;
        RECT 73.725 60.795 73.895 60.965 ;
        RECT 74.185 60.795 74.355 60.965 ;
        RECT 74.645 60.795 74.815 60.965 ;
        RECT 75.105 60.795 75.275 60.965 ;
        RECT 75.565 60.795 75.735 60.965 ;
        RECT 76.025 60.795 76.195 60.965 ;
        RECT 76.485 60.795 76.655 60.965 ;
        RECT 76.945 60.795 77.115 60.965 ;
        RECT 77.405 60.795 77.575 60.965 ;
        RECT 77.865 60.795 78.035 60.965 ;
        RECT 78.325 60.795 78.495 60.965 ;
        RECT 78.785 60.795 78.955 60.965 ;
        RECT 79.245 60.795 79.415 60.965 ;
        RECT 79.705 60.795 79.875 60.965 ;
        RECT 80.165 60.795 80.335 60.965 ;
        RECT 80.625 60.795 80.795 60.965 ;
        RECT 81.085 60.795 81.255 60.965 ;
        RECT 81.545 60.795 81.715 60.965 ;
        RECT 82.005 60.795 82.175 60.965 ;
        RECT 82.465 60.795 82.635 60.965 ;
        RECT 82.925 60.795 83.095 60.965 ;
        RECT 83.385 60.795 83.555 60.965 ;
        RECT 83.845 60.795 84.015 60.965 ;
        RECT 84.305 60.795 84.475 60.965 ;
        RECT 84.765 60.795 84.935 60.965 ;
        RECT 85.225 60.795 85.395 60.965 ;
        RECT 85.685 60.795 85.855 60.965 ;
        RECT 86.145 60.795 86.315 60.965 ;
        RECT 86.605 60.795 86.775 60.965 ;
        RECT 87.065 60.795 87.235 60.965 ;
        RECT 87.525 60.795 87.695 60.965 ;
        RECT 87.985 60.795 88.155 60.965 ;
        RECT 88.445 60.795 88.615 60.965 ;
        RECT 88.905 60.795 89.075 60.965 ;
        RECT 89.365 60.795 89.535 60.965 ;
        RECT 89.825 60.795 89.995 60.965 ;
        RECT 90.285 60.795 90.455 60.965 ;
        RECT 90.745 60.795 90.915 60.965 ;
        RECT 91.205 60.795 91.375 60.965 ;
        RECT 91.665 60.795 91.835 60.965 ;
        RECT 92.125 60.795 92.295 60.965 ;
        RECT 92.585 60.795 92.755 60.965 ;
        RECT 93.045 60.795 93.215 60.965 ;
        RECT 93.505 60.795 93.675 60.965 ;
        RECT 93.965 60.795 94.135 60.965 ;
        RECT 94.425 60.795 94.595 60.965 ;
        RECT 94.885 60.795 95.055 60.965 ;
        RECT 95.345 60.795 95.515 60.965 ;
        RECT 95.805 60.795 95.975 60.965 ;
        RECT 96.265 60.795 96.435 60.965 ;
        RECT 96.725 60.795 96.895 60.965 ;
        RECT 97.185 60.795 97.355 60.965 ;
        RECT 97.645 60.795 97.815 60.965 ;
        RECT 98.105 60.795 98.275 60.965 ;
        RECT 98.565 60.795 98.735 60.965 ;
        RECT 99.025 60.795 99.195 60.965 ;
        RECT 99.485 60.795 99.655 60.965 ;
        RECT 99.945 60.795 100.115 60.965 ;
        RECT 100.405 60.795 100.575 60.965 ;
        RECT 100.865 60.795 101.035 60.965 ;
        RECT 101.325 60.795 101.495 60.965 ;
        RECT 101.785 60.795 101.955 60.965 ;
        RECT 102.245 60.795 102.415 60.965 ;
        RECT 102.705 60.795 102.875 60.965 ;
        RECT 103.165 60.795 103.335 60.965 ;
        RECT 103.625 60.795 103.795 60.965 ;
        RECT 104.085 60.795 104.255 60.965 ;
        RECT 104.545 60.795 104.715 60.965 ;
        RECT 105.005 60.795 105.175 60.965 ;
        RECT 105.465 60.795 105.635 60.965 ;
        RECT 105.925 60.795 106.095 60.965 ;
        RECT 106.385 60.795 106.555 60.965 ;
        RECT 106.845 60.795 107.015 60.965 ;
        RECT 107.305 60.795 107.475 60.965 ;
        RECT 107.765 60.795 107.935 60.965 ;
        RECT 108.225 60.795 108.395 60.965 ;
        RECT 108.685 60.795 108.855 60.965 ;
        RECT 109.145 60.795 109.315 60.965 ;
        RECT 109.605 60.795 109.775 60.965 ;
        RECT 110.065 60.795 110.235 60.965 ;
        RECT 110.525 60.795 110.695 60.965 ;
        RECT 110.985 60.795 111.155 60.965 ;
        RECT 111.445 60.795 111.615 60.965 ;
        RECT 111.905 60.795 112.075 60.965 ;
        RECT 112.365 60.795 112.535 60.965 ;
        RECT 112.825 60.795 112.995 60.965 ;
        RECT 113.285 60.795 113.455 60.965 ;
        RECT 113.745 60.795 113.915 60.965 ;
        RECT 114.205 60.795 114.375 60.965 ;
        RECT 114.665 60.795 114.835 60.965 ;
        RECT 115.125 60.795 115.295 60.965 ;
        RECT 115.585 60.795 115.755 60.965 ;
        RECT 116.045 60.795 116.215 60.965 ;
        RECT 116.505 60.795 116.675 60.965 ;
        RECT 116.965 60.795 117.135 60.965 ;
        RECT 117.425 60.795 117.595 60.965 ;
        RECT 117.885 60.795 118.055 60.965 ;
        RECT 118.345 60.795 118.515 60.965 ;
        RECT 118.805 60.795 118.975 60.965 ;
        RECT 119.265 60.795 119.435 60.965 ;
        RECT 119.725 60.795 119.895 60.965 ;
        RECT 120.185 60.795 120.355 60.965 ;
        RECT 120.645 60.795 120.815 60.965 ;
        RECT 121.105 60.795 121.275 60.965 ;
        RECT 121.565 60.795 121.735 60.965 ;
        RECT 122.025 60.795 122.195 60.965 ;
        RECT 122.485 60.795 122.655 60.965 ;
        RECT 122.945 60.795 123.115 60.965 ;
        RECT 123.405 60.795 123.575 60.965 ;
        RECT 123.865 60.795 124.035 60.965 ;
        RECT 124.325 60.795 124.495 60.965 ;
        RECT 124.785 60.795 124.955 60.965 ;
        RECT 125.245 60.795 125.415 60.965 ;
        RECT 125.705 60.795 125.875 60.965 ;
        RECT 126.165 60.795 126.335 60.965 ;
        RECT 126.625 60.795 126.795 60.965 ;
        RECT 127.085 60.795 127.255 60.965 ;
        RECT 127.545 60.795 127.715 60.965 ;
        RECT 128.005 60.795 128.175 60.965 ;
        RECT 128.465 60.795 128.635 60.965 ;
        RECT 128.925 60.795 129.095 60.965 ;
        RECT 129.385 60.795 129.555 60.965 ;
        RECT 129.845 60.795 130.015 60.965 ;
        RECT 130.305 60.795 130.475 60.965 ;
        RECT 130.765 60.795 130.935 60.965 ;
        RECT 131.225 60.795 131.395 60.965 ;
        RECT 131.685 60.795 131.855 60.965 ;
        RECT 132.145 60.795 132.315 60.965 ;
        RECT 132.605 60.795 132.775 60.965 ;
        RECT 133.065 60.795 133.235 60.965 ;
        RECT 133.525 60.795 133.695 60.965 ;
        RECT 133.985 60.795 134.155 60.965 ;
      LAYER met1 ;
        RECT 45.520 136.800 135.095 137.280 ;
        RECT 45.520 131.360 135.095 131.840 ;
        RECT 45.520 125.920 135.095 126.400 ;
        RECT 45.520 120.480 135.095 120.960 ;
        RECT 45.520 115.040 135.095 115.520 ;
        RECT 45.520 109.600 135.095 110.080 ;
        RECT 45.520 104.160 135.095 104.640 ;
        RECT 45.520 98.720 135.095 99.200 ;
        RECT 45.520 93.280 135.095 93.760 ;
        RECT 45.520 87.840 135.095 88.320 ;
        RECT 45.520 82.400 135.095 82.880 ;
        RECT 45.520 76.960 135.095 77.440 ;
        RECT 45.520 71.520 135.095 72.000 ;
        RECT 45.520 66.080 135.095 66.560 ;
        RECT 45.520 60.640 135.095 61.120 ;
      LAYER via ;
        RECT 66.940 136.910 67.200 137.170 ;
        RECT 67.260 136.910 67.520 137.170 ;
        RECT 67.580 136.910 67.840 137.170 ;
        RECT 67.900 136.910 68.160 137.170 ;
        RECT 68.220 136.910 68.480 137.170 ;
        RECT 89.135 136.910 89.395 137.170 ;
        RECT 89.455 136.910 89.715 137.170 ;
        RECT 89.775 136.910 90.035 137.170 ;
        RECT 90.095 136.910 90.355 137.170 ;
        RECT 90.415 136.910 90.675 137.170 ;
        RECT 111.330 136.910 111.590 137.170 ;
        RECT 111.650 136.910 111.910 137.170 ;
        RECT 111.970 136.910 112.230 137.170 ;
        RECT 112.290 136.910 112.550 137.170 ;
        RECT 112.610 136.910 112.870 137.170 ;
        RECT 133.525 136.910 133.785 137.170 ;
        RECT 133.845 136.910 134.105 137.170 ;
        RECT 134.165 136.910 134.425 137.170 ;
        RECT 134.485 136.910 134.745 137.170 ;
        RECT 134.805 136.910 135.065 137.170 ;
        RECT 66.940 131.470 67.200 131.730 ;
        RECT 67.260 131.470 67.520 131.730 ;
        RECT 67.580 131.470 67.840 131.730 ;
        RECT 67.900 131.470 68.160 131.730 ;
        RECT 68.220 131.470 68.480 131.730 ;
        RECT 89.135 131.470 89.395 131.730 ;
        RECT 89.455 131.470 89.715 131.730 ;
        RECT 89.775 131.470 90.035 131.730 ;
        RECT 90.095 131.470 90.355 131.730 ;
        RECT 90.415 131.470 90.675 131.730 ;
        RECT 111.330 131.470 111.590 131.730 ;
        RECT 111.650 131.470 111.910 131.730 ;
        RECT 111.970 131.470 112.230 131.730 ;
        RECT 112.290 131.470 112.550 131.730 ;
        RECT 112.610 131.470 112.870 131.730 ;
        RECT 133.525 131.470 133.785 131.730 ;
        RECT 133.845 131.470 134.105 131.730 ;
        RECT 134.165 131.470 134.425 131.730 ;
        RECT 134.485 131.470 134.745 131.730 ;
        RECT 134.805 131.470 135.065 131.730 ;
        RECT 66.940 126.030 67.200 126.290 ;
        RECT 67.260 126.030 67.520 126.290 ;
        RECT 67.580 126.030 67.840 126.290 ;
        RECT 67.900 126.030 68.160 126.290 ;
        RECT 68.220 126.030 68.480 126.290 ;
        RECT 89.135 126.030 89.395 126.290 ;
        RECT 89.455 126.030 89.715 126.290 ;
        RECT 89.775 126.030 90.035 126.290 ;
        RECT 90.095 126.030 90.355 126.290 ;
        RECT 90.415 126.030 90.675 126.290 ;
        RECT 111.330 126.030 111.590 126.290 ;
        RECT 111.650 126.030 111.910 126.290 ;
        RECT 111.970 126.030 112.230 126.290 ;
        RECT 112.290 126.030 112.550 126.290 ;
        RECT 112.610 126.030 112.870 126.290 ;
        RECT 133.525 126.030 133.785 126.290 ;
        RECT 133.845 126.030 134.105 126.290 ;
        RECT 134.165 126.030 134.425 126.290 ;
        RECT 134.485 126.030 134.745 126.290 ;
        RECT 134.805 126.030 135.065 126.290 ;
        RECT 66.940 120.590 67.200 120.850 ;
        RECT 67.260 120.590 67.520 120.850 ;
        RECT 67.580 120.590 67.840 120.850 ;
        RECT 67.900 120.590 68.160 120.850 ;
        RECT 68.220 120.590 68.480 120.850 ;
        RECT 89.135 120.590 89.395 120.850 ;
        RECT 89.455 120.590 89.715 120.850 ;
        RECT 89.775 120.590 90.035 120.850 ;
        RECT 90.095 120.590 90.355 120.850 ;
        RECT 90.415 120.590 90.675 120.850 ;
        RECT 111.330 120.590 111.590 120.850 ;
        RECT 111.650 120.590 111.910 120.850 ;
        RECT 111.970 120.590 112.230 120.850 ;
        RECT 112.290 120.590 112.550 120.850 ;
        RECT 112.610 120.590 112.870 120.850 ;
        RECT 133.525 120.590 133.785 120.850 ;
        RECT 133.845 120.590 134.105 120.850 ;
        RECT 134.165 120.590 134.425 120.850 ;
        RECT 134.485 120.590 134.745 120.850 ;
        RECT 134.805 120.590 135.065 120.850 ;
        RECT 66.940 115.150 67.200 115.410 ;
        RECT 67.260 115.150 67.520 115.410 ;
        RECT 67.580 115.150 67.840 115.410 ;
        RECT 67.900 115.150 68.160 115.410 ;
        RECT 68.220 115.150 68.480 115.410 ;
        RECT 89.135 115.150 89.395 115.410 ;
        RECT 89.455 115.150 89.715 115.410 ;
        RECT 89.775 115.150 90.035 115.410 ;
        RECT 90.095 115.150 90.355 115.410 ;
        RECT 90.415 115.150 90.675 115.410 ;
        RECT 111.330 115.150 111.590 115.410 ;
        RECT 111.650 115.150 111.910 115.410 ;
        RECT 111.970 115.150 112.230 115.410 ;
        RECT 112.290 115.150 112.550 115.410 ;
        RECT 112.610 115.150 112.870 115.410 ;
        RECT 133.525 115.150 133.785 115.410 ;
        RECT 133.845 115.150 134.105 115.410 ;
        RECT 134.165 115.150 134.425 115.410 ;
        RECT 134.485 115.150 134.745 115.410 ;
        RECT 134.805 115.150 135.065 115.410 ;
        RECT 66.940 109.710 67.200 109.970 ;
        RECT 67.260 109.710 67.520 109.970 ;
        RECT 67.580 109.710 67.840 109.970 ;
        RECT 67.900 109.710 68.160 109.970 ;
        RECT 68.220 109.710 68.480 109.970 ;
        RECT 89.135 109.710 89.395 109.970 ;
        RECT 89.455 109.710 89.715 109.970 ;
        RECT 89.775 109.710 90.035 109.970 ;
        RECT 90.095 109.710 90.355 109.970 ;
        RECT 90.415 109.710 90.675 109.970 ;
        RECT 111.330 109.710 111.590 109.970 ;
        RECT 111.650 109.710 111.910 109.970 ;
        RECT 111.970 109.710 112.230 109.970 ;
        RECT 112.290 109.710 112.550 109.970 ;
        RECT 112.610 109.710 112.870 109.970 ;
        RECT 133.525 109.710 133.785 109.970 ;
        RECT 133.845 109.710 134.105 109.970 ;
        RECT 134.165 109.710 134.425 109.970 ;
        RECT 134.485 109.710 134.745 109.970 ;
        RECT 134.805 109.710 135.065 109.970 ;
        RECT 66.940 104.270 67.200 104.530 ;
        RECT 67.260 104.270 67.520 104.530 ;
        RECT 67.580 104.270 67.840 104.530 ;
        RECT 67.900 104.270 68.160 104.530 ;
        RECT 68.220 104.270 68.480 104.530 ;
        RECT 89.135 104.270 89.395 104.530 ;
        RECT 89.455 104.270 89.715 104.530 ;
        RECT 89.775 104.270 90.035 104.530 ;
        RECT 90.095 104.270 90.355 104.530 ;
        RECT 90.415 104.270 90.675 104.530 ;
        RECT 111.330 104.270 111.590 104.530 ;
        RECT 111.650 104.270 111.910 104.530 ;
        RECT 111.970 104.270 112.230 104.530 ;
        RECT 112.290 104.270 112.550 104.530 ;
        RECT 112.610 104.270 112.870 104.530 ;
        RECT 133.525 104.270 133.785 104.530 ;
        RECT 133.845 104.270 134.105 104.530 ;
        RECT 134.165 104.270 134.425 104.530 ;
        RECT 134.485 104.270 134.745 104.530 ;
        RECT 134.805 104.270 135.065 104.530 ;
        RECT 66.940 98.830 67.200 99.090 ;
        RECT 67.260 98.830 67.520 99.090 ;
        RECT 67.580 98.830 67.840 99.090 ;
        RECT 67.900 98.830 68.160 99.090 ;
        RECT 68.220 98.830 68.480 99.090 ;
        RECT 89.135 98.830 89.395 99.090 ;
        RECT 89.455 98.830 89.715 99.090 ;
        RECT 89.775 98.830 90.035 99.090 ;
        RECT 90.095 98.830 90.355 99.090 ;
        RECT 90.415 98.830 90.675 99.090 ;
        RECT 111.330 98.830 111.590 99.090 ;
        RECT 111.650 98.830 111.910 99.090 ;
        RECT 111.970 98.830 112.230 99.090 ;
        RECT 112.290 98.830 112.550 99.090 ;
        RECT 112.610 98.830 112.870 99.090 ;
        RECT 133.525 98.830 133.785 99.090 ;
        RECT 133.845 98.830 134.105 99.090 ;
        RECT 134.165 98.830 134.425 99.090 ;
        RECT 134.485 98.830 134.745 99.090 ;
        RECT 134.805 98.830 135.065 99.090 ;
        RECT 66.940 93.390 67.200 93.650 ;
        RECT 67.260 93.390 67.520 93.650 ;
        RECT 67.580 93.390 67.840 93.650 ;
        RECT 67.900 93.390 68.160 93.650 ;
        RECT 68.220 93.390 68.480 93.650 ;
        RECT 89.135 93.390 89.395 93.650 ;
        RECT 89.455 93.390 89.715 93.650 ;
        RECT 89.775 93.390 90.035 93.650 ;
        RECT 90.095 93.390 90.355 93.650 ;
        RECT 90.415 93.390 90.675 93.650 ;
        RECT 111.330 93.390 111.590 93.650 ;
        RECT 111.650 93.390 111.910 93.650 ;
        RECT 111.970 93.390 112.230 93.650 ;
        RECT 112.290 93.390 112.550 93.650 ;
        RECT 112.610 93.390 112.870 93.650 ;
        RECT 133.525 93.390 133.785 93.650 ;
        RECT 133.845 93.390 134.105 93.650 ;
        RECT 134.165 93.390 134.425 93.650 ;
        RECT 134.485 93.390 134.745 93.650 ;
        RECT 134.805 93.390 135.065 93.650 ;
        RECT 66.940 87.950 67.200 88.210 ;
        RECT 67.260 87.950 67.520 88.210 ;
        RECT 67.580 87.950 67.840 88.210 ;
        RECT 67.900 87.950 68.160 88.210 ;
        RECT 68.220 87.950 68.480 88.210 ;
        RECT 89.135 87.950 89.395 88.210 ;
        RECT 89.455 87.950 89.715 88.210 ;
        RECT 89.775 87.950 90.035 88.210 ;
        RECT 90.095 87.950 90.355 88.210 ;
        RECT 90.415 87.950 90.675 88.210 ;
        RECT 111.330 87.950 111.590 88.210 ;
        RECT 111.650 87.950 111.910 88.210 ;
        RECT 111.970 87.950 112.230 88.210 ;
        RECT 112.290 87.950 112.550 88.210 ;
        RECT 112.610 87.950 112.870 88.210 ;
        RECT 133.525 87.950 133.785 88.210 ;
        RECT 133.845 87.950 134.105 88.210 ;
        RECT 134.165 87.950 134.425 88.210 ;
        RECT 134.485 87.950 134.745 88.210 ;
        RECT 134.805 87.950 135.065 88.210 ;
        RECT 66.940 82.510 67.200 82.770 ;
        RECT 67.260 82.510 67.520 82.770 ;
        RECT 67.580 82.510 67.840 82.770 ;
        RECT 67.900 82.510 68.160 82.770 ;
        RECT 68.220 82.510 68.480 82.770 ;
        RECT 89.135 82.510 89.395 82.770 ;
        RECT 89.455 82.510 89.715 82.770 ;
        RECT 89.775 82.510 90.035 82.770 ;
        RECT 90.095 82.510 90.355 82.770 ;
        RECT 90.415 82.510 90.675 82.770 ;
        RECT 111.330 82.510 111.590 82.770 ;
        RECT 111.650 82.510 111.910 82.770 ;
        RECT 111.970 82.510 112.230 82.770 ;
        RECT 112.290 82.510 112.550 82.770 ;
        RECT 112.610 82.510 112.870 82.770 ;
        RECT 133.525 82.510 133.785 82.770 ;
        RECT 133.845 82.510 134.105 82.770 ;
        RECT 134.165 82.510 134.425 82.770 ;
        RECT 134.485 82.510 134.745 82.770 ;
        RECT 134.805 82.510 135.065 82.770 ;
        RECT 66.940 77.070 67.200 77.330 ;
        RECT 67.260 77.070 67.520 77.330 ;
        RECT 67.580 77.070 67.840 77.330 ;
        RECT 67.900 77.070 68.160 77.330 ;
        RECT 68.220 77.070 68.480 77.330 ;
        RECT 89.135 77.070 89.395 77.330 ;
        RECT 89.455 77.070 89.715 77.330 ;
        RECT 89.775 77.070 90.035 77.330 ;
        RECT 90.095 77.070 90.355 77.330 ;
        RECT 90.415 77.070 90.675 77.330 ;
        RECT 111.330 77.070 111.590 77.330 ;
        RECT 111.650 77.070 111.910 77.330 ;
        RECT 111.970 77.070 112.230 77.330 ;
        RECT 112.290 77.070 112.550 77.330 ;
        RECT 112.610 77.070 112.870 77.330 ;
        RECT 133.525 77.070 133.785 77.330 ;
        RECT 133.845 77.070 134.105 77.330 ;
        RECT 134.165 77.070 134.425 77.330 ;
        RECT 134.485 77.070 134.745 77.330 ;
        RECT 134.805 77.070 135.065 77.330 ;
        RECT 66.940 71.630 67.200 71.890 ;
        RECT 67.260 71.630 67.520 71.890 ;
        RECT 67.580 71.630 67.840 71.890 ;
        RECT 67.900 71.630 68.160 71.890 ;
        RECT 68.220 71.630 68.480 71.890 ;
        RECT 89.135 71.630 89.395 71.890 ;
        RECT 89.455 71.630 89.715 71.890 ;
        RECT 89.775 71.630 90.035 71.890 ;
        RECT 90.095 71.630 90.355 71.890 ;
        RECT 90.415 71.630 90.675 71.890 ;
        RECT 111.330 71.630 111.590 71.890 ;
        RECT 111.650 71.630 111.910 71.890 ;
        RECT 111.970 71.630 112.230 71.890 ;
        RECT 112.290 71.630 112.550 71.890 ;
        RECT 112.610 71.630 112.870 71.890 ;
        RECT 133.525 71.630 133.785 71.890 ;
        RECT 133.845 71.630 134.105 71.890 ;
        RECT 134.165 71.630 134.425 71.890 ;
        RECT 134.485 71.630 134.745 71.890 ;
        RECT 134.805 71.630 135.065 71.890 ;
        RECT 66.940 66.190 67.200 66.450 ;
        RECT 67.260 66.190 67.520 66.450 ;
        RECT 67.580 66.190 67.840 66.450 ;
        RECT 67.900 66.190 68.160 66.450 ;
        RECT 68.220 66.190 68.480 66.450 ;
        RECT 89.135 66.190 89.395 66.450 ;
        RECT 89.455 66.190 89.715 66.450 ;
        RECT 89.775 66.190 90.035 66.450 ;
        RECT 90.095 66.190 90.355 66.450 ;
        RECT 90.415 66.190 90.675 66.450 ;
        RECT 111.330 66.190 111.590 66.450 ;
        RECT 111.650 66.190 111.910 66.450 ;
        RECT 111.970 66.190 112.230 66.450 ;
        RECT 112.290 66.190 112.550 66.450 ;
        RECT 112.610 66.190 112.870 66.450 ;
        RECT 133.525 66.190 133.785 66.450 ;
        RECT 133.845 66.190 134.105 66.450 ;
        RECT 134.165 66.190 134.425 66.450 ;
        RECT 134.485 66.190 134.745 66.450 ;
        RECT 134.805 66.190 135.065 66.450 ;
        RECT 66.940 60.750 67.200 61.010 ;
        RECT 67.260 60.750 67.520 61.010 ;
        RECT 67.580 60.750 67.840 61.010 ;
        RECT 67.900 60.750 68.160 61.010 ;
        RECT 68.220 60.750 68.480 61.010 ;
        RECT 89.135 60.750 89.395 61.010 ;
        RECT 89.455 60.750 89.715 61.010 ;
        RECT 89.775 60.750 90.035 61.010 ;
        RECT 90.095 60.750 90.355 61.010 ;
        RECT 90.415 60.750 90.675 61.010 ;
        RECT 111.330 60.750 111.590 61.010 ;
        RECT 111.650 60.750 111.910 61.010 ;
        RECT 111.970 60.750 112.230 61.010 ;
        RECT 112.290 60.750 112.550 61.010 ;
        RECT 112.610 60.750 112.870 61.010 ;
        RECT 133.525 60.750 133.785 61.010 ;
        RECT 133.845 60.750 134.105 61.010 ;
        RECT 134.165 60.750 134.425 61.010 ;
        RECT 134.485 60.750 134.745 61.010 ;
        RECT 134.805 60.750 135.065 61.010 ;
      LAYER met2 ;
        RECT 66.940 136.855 68.480 137.225 ;
        RECT 89.135 136.855 90.675 137.225 ;
        RECT 111.330 136.855 112.870 137.225 ;
        RECT 133.525 136.855 135.065 137.225 ;
        RECT 66.940 131.415 68.480 131.785 ;
        RECT 89.135 131.415 90.675 131.785 ;
        RECT 111.330 131.415 112.870 131.785 ;
        RECT 133.525 131.415 135.065 131.785 ;
        RECT 66.940 125.975 68.480 126.345 ;
        RECT 89.135 125.975 90.675 126.345 ;
        RECT 111.330 125.975 112.870 126.345 ;
        RECT 133.525 125.975 135.065 126.345 ;
        RECT 66.940 120.535 68.480 120.905 ;
        RECT 89.135 120.535 90.675 120.905 ;
        RECT 111.330 120.535 112.870 120.905 ;
        RECT 133.525 120.535 135.065 120.905 ;
        RECT 66.940 115.095 68.480 115.465 ;
        RECT 89.135 115.095 90.675 115.465 ;
        RECT 111.330 115.095 112.870 115.465 ;
        RECT 133.525 115.095 135.065 115.465 ;
        RECT 66.940 109.655 68.480 110.025 ;
        RECT 89.135 109.655 90.675 110.025 ;
        RECT 111.330 109.655 112.870 110.025 ;
        RECT 133.525 109.655 135.065 110.025 ;
        RECT 66.940 104.215 68.480 104.585 ;
        RECT 89.135 104.215 90.675 104.585 ;
        RECT 111.330 104.215 112.870 104.585 ;
        RECT 133.525 104.215 135.065 104.585 ;
        RECT 66.940 98.775 68.480 99.145 ;
        RECT 89.135 98.775 90.675 99.145 ;
        RECT 111.330 98.775 112.870 99.145 ;
        RECT 133.525 98.775 135.065 99.145 ;
        RECT 66.940 93.335 68.480 93.705 ;
        RECT 89.135 93.335 90.675 93.705 ;
        RECT 111.330 93.335 112.870 93.705 ;
        RECT 133.525 93.335 135.065 93.705 ;
        RECT 66.940 87.895 68.480 88.265 ;
        RECT 89.135 87.895 90.675 88.265 ;
        RECT 111.330 87.895 112.870 88.265 ;
        RECT 133.525 87.895 135.065 88.265 ;
        RECT 66.940 82.455 68.480 82.825 ;
        RECT 89.135 82.455 90.675 82.825 ;
        RECT 111.330 82.455 112.870 82.825 ;
        RECT 133.525 82.455 135.065 82.825 ;
        RECT 66.940 77.015 68.480 77.385 ;
        RECT 89.135 77.015 90.675 77.385 ;
        RECT 111.330 77.015 112.870 77.385 ;
        RECT 133.525 77.015 135.065 77.385 ;
        RECT 66.940 71.575 68.480 71.945 ;
        RECT 89.135 71.575 90.675 71.945 ;
        RECT 111.330 71.575 112.870 71.945 ;
        RECT 133.525 71.575 135.065 71.945 ;
        RECT 66.940 66.135 68.480 66.505 ;
        RECT 89.135 66.135 90.675 66.505 ;
        RECT 111.330 66.135 112.870 66.505 ;
        RECT 133.525 66.135 135.065 66.505 ;
        RECT 66.940 60.695 68.480 61.065 ;
        RECT 89.135 60.695 90.675 61.065 ;
        RECT 111.330 60.695 112.870 61.065 ;
        RECT 133.525 60.695 135.065 61.065 ;
      LAYER via2 ;
        RECT 66.970 136.900 67.250 137.180 ;
        RECT 67.370 136.900 67.650 137.180 ;
        RECT 67.770 136.900 68.050 137.180 ;
        RECT 68.170 136.900 68.450 137.180 ;
        RECT 89.165 136.900 89.445 137.180 ;
        RECT 89.565 136.900 89.845 137.180 ;
        RECT 89.965 136.900 90.245 137.180 ;
        RECT 90.365 136.900 90.645 137.180 ;
        RECT 111.360 136.900 111.640 137.180 ;
        RECT 111.760 136.900 112.040 137.180 ;
        RECT 112.160 136.900 112.440 137.180 ;
        RECT 112.560 136.900 112.840 137.180 ;
        RECT 133.555 136.900 133.835 137.180 ;
        RECT 133.955 136.900 134.235 137.180 ;
        RECT 134.355 136.900 134.635 137.180 ;
        RECT 134.755 136.900 135.035 137.180 ;
        RECT 66.970 131.460 67.250 131.740 ;
        RECT 67.370 131.460 67.650 131.740 ;
        RECT 67.770 131.460 68.050 131.740 ;
        RECT 68.170 131.460 68.450 131.740 ;
        RECT 89.165 131.460 89.445 131.740 ;
        RECT 89.565 131.460 89.845 131.740 ;
        RECT 89.965 131.460 90.245 131.740 ;
        RECT 90.365 131.460 90.645 131.740 ;
        RECT 111.360 131.460 111.640 131.740 ;
        RECT 111.760 131.460 112.040 131.740 ;
        RECT 112.160 131.460 112.440 131.740 ;
        RECT 112.560 131.460 112.840 131.740 ;
        RECT 133.555 131.460 133.835 131.740 ;
        RECT 133.955 131.460 134.235 131.740 ;
        RECT 134.355 131.460 134.635 131.740 ;
        RECT 134.755 131.460 135.035 131.740 ;
        RECT 66.970 126.020 67.250 126.300 ;
        RECT 67.370 126.020 67.650 126.300 ;
        RECT 67.770 126.020 68.050 126.300 ;
        RECT 68.170 126.020 68.450 126.300 ;
        RECT 89.165 126.020 89.445 126.300 ;
        RECT 89.565 126.020 89.845 126.300 ;
        RECT 89.965 126.020 90.245 126.300 ;
        RECT 90.365 126.020 90.645 126.300 ;
        RECT 111.360 126.020 111.640 126.300 ;
        RECT 111.760 126.020 112.040 126.300 ;
        RECT 112.160 126.020 112.440 126.300 ;
        RECT 112.560 126.020 112.840 126.300 ;
        RECT 133.555 126.020 133.835 126.300 ;
        RECT 133.955 126.020 134.235 126.300 ;
        RECT 134.355 126.020 134.635 126.300 ;
        RECT 134.755 126.020 135.035 126.300 ;
        RECT 66.970 120.580 67.250 120.860 ;
        RECT 67.370 120.580 67.650 120.860 ;
        RECT 67.770 120.580 68.050 120.860 ;
        RECT 68.170 120.580 68.450 120.860 ;
        RECT 89.165 120.580 89.445 120.860 ;
        RECT 89.565 120.580 89.845 120.860 ;
        RECT 89.965 120.580 90.245 120.860 ;
        RECT 90.365 120.580 90.645 120.860 ;
        RECT 111.360 120.580 111.640 120.860 ;
        RECT 111.760 120.580 112.040 120.860 ;
        RECT 112.160 120.580 112.440 120.860 ;
        RECT 112.560 120.580 112.840 120.860 ;
        RECT 133.555 120.580 133.835 120.860 ;
        RECT 133.955 120.580 134.235 120.860 ;
        RECT 134.355 120.580 134.635 120.860 ;
        RECT 134.755 120.580 135.035 120.860 ;
        RECT 66.970 115.140 67.250 115.420 ;
        RECT 67.370 115.140 67.650 115.420 ;
        RECT 67.770 115.140 68.050 115.420 ;
        RECT 68.170 115.140 68.450 115.420 ;
        RECT 89.165 115.140 89.445 115.420 ;
        RECT 89.565 115.140 89.845 115.420 ;
        RECT 89.965 115.140 90.245 115.420 ;
        RECT 90.365 115.140 90.645 115.420 ;
        RECT 111.360 115.140 111.640 115.420 ;
        RECT 111.760 115.140 112.040 115.420 ;
        RECT 112.160 115.140 112.440 115.420 ;
        RECT 112.560 115.140 112.840 115.420 ;
        RECT 133.555 115.140 133.835 115.420 ;
        RECT 133.955 115.140 134.235 115.420 ;
        RECT 134.355 115.140 134.635 115.420 ;
        RECT 134.755 115.140 135.035 115.420 ;
        RECT 66.970 109.700 67.250 109.980 ;
        RECT 67.370 109.700 67.650 109.980 ;
        RECT 67.770 109.700 68.050 109.980 ;
        RECT 68.170 109.700 68.450 109.980 ;
        RECT 89.165 109.700 89.445 109.980 ;
        RECT 89.565 109.700 89.845 109.980 ;
        RECT 89.965 109.700 90.245 109.980 ;
        RECT 90.365 109.700 90.645 109.980 ;
        RECT 111.360 109.700 111.640 109.980 ;
        RECT 111.760 109.700 112.040 109.980 ;
        RECT 112.160 109.700 112.440 109.980 ;
        RECT 112.560 109.700 112.840 109.980 ;
        RECT 133.555 109.700 133.835 109.980 ;
        RECT 133.955 109.700 134.235 109.980 ;
        RECT 134.355 109.700 134.635 109.980 ;
        RECT 134.755 109.700 135.035 109.980 ;
        RECT 66.970 104.260 67.250 104.540 ;
        RECT 67.370 104.260 67.650 104.540 ;
        RECT 67.770 104.260 68.050 104.540 ;
        RECT 68.170 104.260 68.450 104.540 ;
        RECT 89.165 104.260 89.445 104.540 ;
        RECT 89.565 104.260 89.845 104.540 ;
        RECT 89.965 104.260 90.245 104.540 ;
        RECT 90.365 104.260 90.645 104.540 ;
        RECT 111.360 104.260 111.640 104.540 ;
        RECT 111.760 104.260 112.040 104.540 ;
        RECT 112.160 104.260 112.440 104.540 ;
        RECT 112.560 104.260 112.840 104.540 ;
        RECT 133.555 104.260 133.835 104.540 ;
        RECT 133.955 104.260 134.235 104.540 ;
        RECT 134.355 104.260 134.635 104.540 ;
        RECT 134.755 104.260 135.035 104.540 ;
        RECT 66.970 98.820 67.250 99.100 ;
        RECT 67.370 98.820 67.650 99.100 ;
        RECT 67.770 98.820 68.050 99.100 ;
        RECT 68.170 98.820 68.450 99.100 ;
        RECT 89.165 98.820 89.445 99.100 ;
        RECT 89.565 98.820 89.845 99.100 ;
        RECT 89.965 98.820 90.245 99.100 ;
        RECT 90.365 98.820 90.645 99.100 ;
        RECT 111.360 98.820 111.640 99.100 ;
        RECT 111.760 98.820 112.040 99.100 ;
        RECT 112.160 98.820 112.440 99.100 ;
        RECT 112.560 98.820 112.840 99.100 ;
        RECT 133.555 98.820 133.835 99.100 ;
        RECT 133.955 98.820 134.235 99.100 ;
        RECT 134.355 98.820 134.635 99.100 ;
        RECT 134.755 98.820 135.035 99.100 ;
        RECT 66.970 93.380 67.250 93.660 ;
        RECT 67.370 93.380 67.650 93.660 ;
        RECT 67.770 93.380 68.050 93.660 ;
        RECT 68.170 93.380 68.450 93.660 ;
        RECT 89.165 93.380 89.445 93.660 ;
        RECT 89.565 93.380 89.845 93.660 ;
        RECT 89.965 93.380 90.245 93.660 ;
        RECT 90.365 93.380 90.645 93.660 ;
        RECT 111.360 93.380 111.640 93.660 ;
        RECT 111.760 93.380 112.040 93.660 ;
        RECT 112.160 93.380 112.440 93.660 ;
        RECT 112.560 93.380 112.840 93.660 ;
        RECT 133.555 93.380 133.835 93.660 ;
        RECT 133.955 93.380 134.235 93.660 ;
        RECT 134.355 93.380 134.635 93.660 ;
        RECT 134.755 93.380 135.035 93.660 ;
        RECT 66.970 87.940 67.250 88.220 ;
        RECT 67.370 87.940 67.650 88.220 ;
        RECT 67.770 87.940 68.050 88.220 ;
        RECT 68.170 87.940 68.450 88.220 ;
        RECT 89.165 87.940 89.445 88.220 ;
        RECT 89.565 87.940 89.845 88.220 ;
        RECT 89.965 87.940 90.245 88.220 ;
        RECT 90.365 87.940 90.645 88.220 ;
        RECT 111.360 87.940 111.640 88.220 ;
        RECT 111.760 87.940 112.040 88.220 ;
        RECT 112.160 87.940 112.440 88.220 ;
        RECT 112.560 87.940 112.840 88.220 ;
        RECT 133.555 87.940 133.835 88.220 ;
        RECT 133.955 87.940 134.235 88.220 ;
        RECT 134.355 87.940 134.635 88.220 ;
        RECT 134.755 87.940 135.035 88.220 ;
        RECT 66.970 82.500 67.250 82.780 ;
        RECT 67.370 82.500 67.650 82.780 ;
        RECT 67.770 82.500 68.050 82.780 ;
        RECT 68.170 82.500 68.450 82.780 ;
        RECT 89.165 82.500 89.445 82.780 ;
        RECT 89.565 82.500 89.845 82.780 ;
        RECT 89.965 82.500 90.245 82.780 ;
        RECT 90.365 82.500 90.645 82.780 ;
        RECT 111.360 82.500 111.640 82.780 ;
        RECT 111.760 82.500 112.040 82.780 ;
        RECT 112.160 82.500 112.440 82.780 ;
        RECT 112.560 82.500 112.840 82.780 ;
        RECT 133.555 82.500 133.835 82.780 ;
        RECT 133.955 82.500 134.235 82.780 ;
        RECT 134.355 82.500 134.635 82.780 ;
        RECT 134.755 82.500 135.035 82.780 ;
        RECT 66.970 77.060 67.250 77.340 ;
        RECT 67.370 77.060 67.650 77.340 ;
        RECT 67.770 77.060 68.050 77.340 ;
        RECT 68.170 77.060 68.450 77.340 ;
        RECT 89.165 77.060 89.445 77.340 ;
        RECT 89.565 77.060 89.845 77.340 ;
        RECT 89.965 77.060 90.245 77.340 ;
        RECT 90.365 77.060 90.645 77.340 ;
        RECT 111.360 77.060 111.640 77.340 ;
        RECT 111.760 77.060 112.040 77.340 ;
        RECT 112.160 77.060 112.440 77.340 ;
        RECT 112.560 77.060 112.840 77.340 ;
        RECT 133.555 77.060 133.835 77.340 ;
        RECT 133.955 77.060 134.235 77.340 ;
        RECT 134.355 77.060 134.635 77.340 ;
        RECT 134.755 77.060 135.035 77.340 ;
        RECT 66.970 71.620 67.250 71.900 ;
        RECT 67.370 71.620 67.650 71.900 ;
        RECT 67.770 71.620 68.050 71.900 ;
        RECT 68.170 71.620 68.450 71.900 ;
        RECT 89.165 71.620 89.445 71.900 ;
        RECT 89.565 71.620 89.845 71.900 ;
        RECT 89.965 71.620 90.245 71.900 ;
        RECT 90.365 71.620 90.645 71.900 ;
        RECT 111.360 71.620 111.640 71.900 ;
        RECT 111.760 71.620 112.040 71.900 ;
        RECT 112.160 71.620 112.440 71.900 ;
        RECT 112.560 71.620 112.840 71.900 ;
        RECT 133.555 71.620 133.835 71.900 ;
        RECT 133.955 71.620 134.235 71.900 ;
        RECT 134.355 71.620 134.635 71.900 ;
        RECT 134.755 71.620 135.035 71.900 ;
        RECT 66.970 66.180 67.250 66.460 ;
        RECT 67.370 66.180 67.650 66.460 ;
        RECT 67.770 66.180 68.050 66.460 ;
        RECT 68.170 66.180 68.450 66.460 ;
        RECT 89.165 66.180 89.445 66.460 ;
        RECT 89.565 66.180 89.845 66.460 ;
        RECT 89.965 66.180 90.245 66.460 ;
        RECT 90.365 66.180 90.645 66.460 ;
        RECT 111.360 66.180 111.640 66.460 ;
        RECT 111.760 66.180 112.040 66.460 ;
        RECT 112.160 66.180 112.440 66.460 ;
        RECT 112.560 66.180 112.840 66.460 ;
        RECT 133.555 66.180 133.835 66.460 ;
        RECT 133.955 66.180 134.235 66.460 ;
        RECT 134.355 66.180 134.635 66.460 ;
        RECT 134.755 66.180 135.035 66.460 ;
        RECT 66.970 60.740 67.250 61.020 ;
        RECT 67.370 60.740 67.650 61.020 ;
        RECT 67.770 60.740 68.050 61.020 ;
        RECT 68.170 60.740 68.450 61.020 ;
        RECT 89.165 60.740 89.445 61.020 ;
        RECT 89.565 60.740 89.845 61.020 ;
        RECT 89.965 60.740 90.245 61.020 ;
        RECT 90.365 60.740 90.645 61.020 ;
        RECT 111.360 60.740 111.640 61.020 ;
        RECT 111.760 60.740 112.040 61.020 ;
        RECT 112.160 60.740 112.440 61.020 ;
        RECT 112.560 60.740 112.840 61.020 ;
        RECT 133.555 60.740 133.835 61.020 ;
        RECT 133.955 60.740 134.235 61.020 ;
        RECT 134.355 60.740 134.635 61.020 ;
        RECT 134.755 60.740 135.035 61.020 ;
      LAYER met3 ;
        RECT 66.920 136.875 68.500 137.205 ;
        RECT 89.115 136.875 90.695 137.205 ;
        RECT 111.310 136.875 112.890 137.205 ;
        RECT 133.505 136.875 135.085 137.205 ;
        RECT 66.920 131.435 68.500 131.765 ;
        RECT 89.115 131.435 90.695 131.765 ;
        RECT 111.310 131.435 112.890 131.765 ;
        RECT 133.505 131.435 135.085 131.765 ;
        RECT 66.920 125.995 68.500 126.325 ;
        RECT 89.115 125.995 90.695 126.325 ;
        RECT 111.310 125.995 112.890 126.325 ;
        RECT 133.505 125.995 135.085 126.325 ;
        RECT 66.920 120.555 68.500 120.885 ;
        RECT 89.115 120.555 90.695 120.885 ;
        RECT 111.310 120.555 112.890 120.885 ;
        RECT 133.505 120.555 135.085 120.885 ;
        RECT 66.920 115.115 68.500 115.445 ;
        RECT 89.115 115.115 90.695 115.445 ;
        RECT 111.310 115.115 112.890 115.445 ;
        RECT 133.505 115.115 135.085 115.445 ;
        RECT 66.920 109.675 68.500 110.005 ;
        RECT 89.115 109.675 90.695 110.005 ;
        RECT 111.310 109.675 112.890 110.005 ;
        RECT 133.505 109.675 135.085 110.005 ;
        RECT 66.920 104.235 68.500 104.565 ;
        RECT 89.115 104.235 90.695 104.565 ;
        RECT 111.310 104.235 112.890 104.565 ;
        RECT 133.505 104.235 135.085 104.565 ;
        RECT 66.920 98.795 68.500 99.125 ;
        RECT 89.115 98.795 90.695 99.125 ;
        RECT 111.310 98.795 112.890 99.125 ;
        RECT 133.505 98.795 135.085 99.125 ;
        RECT 66.920 93.355 68.500 93.685 ;
        RECT 89.115 93.355 90.695 93.685 ;
        RECT 111.310 93.355 112.890 93.685 ;
        RECT 133.505 93.355 135.085 93.685 ;
        RECT 66.920 87.915 68.500 88.245 ;
        RECT 89.115 87.915 90.695 88.245 ;
        RECT 111.310 87.915 112.890 88.245 ;
        RECT 133.505 87.915 135.085 88.245 ;
        RECT 66.920 82.475 68.500 82.805 ;
        RECT 89.115 82.475 90.695 82.805 ;
        RECT 111.310 82.475 112.890 82.805 ;
        RECT 133.505 82.475 135.085 82.805 ;
        RECT 66.920 77.035 68.500 77.365 ;
        RECT 89.115 77.035 90.695 77.365 ;
        RECT 111.310 77.035 112.890 77.365 ;
        RECT 133.505 77.035 135.085 77.365 ;
        RECT 66.920 71.595 68.500 71.925 ;
        RECT 89.115 71.595 90.695 71.925 ;
        RECT 111.310 71.595 112.890 71.925 ;
        RECT 133.505 71.595 135.085 71.925 ;
        RECT 66.920 66.155 68.500 66.485 ;
        RECT 89.115 66.155 90.695 66.485 ;
        RECT 111.310 66.155 112.890 66.485 ;
        RECT 133.505 66.155 135.085 66.485 ;
        RECT 66.920 60.715 68.500 61.045 ;
        RECT 89.115 60.715 90.695 61.045 ;
        RECT 111.310 60.715 112.890 61.045 ;
        RECT 133.505 60.715 135.085 61.045 ;
      LAYER via3 ;
        RECT 66.950 136.880 67.270 137.200 ;
        RECT 67.350 136.880 67.670 137.200 ;
        RECT 67.750 136.880 68.070 137.200 ;
        RECT 68.150 136.880 68.470 137.200 ;
        RECT 89.145 136.880 89.465 137.200 ;
        RECT 89.545 136.880 89.865 137.200 ;
        RECT 89.945 136.880 90.265 137.200 ;
        RECT 90.345 136.880 90.665 137.200 ;
        RECT 111.340 136.880 111.660 137.200 ;
        RECT 111.740 136.880 112.060 137.200 ;
        RECT 112.140 136.880 112.460 137.200 ;
        RECT 112.540 136.880 112.860 137.200 ;
        RECT 133.535 136.880 133.855 137.200 ;
        RECT 133.935 136.880 134.255 137.200 ;
        RECT 134.335 136.880 134.655 137.200 ;
        RECT 134.735 136.880 135.055 137.200 ;
        RECT 66.950 131.440 67.270 131.760 ;
        RECT 67.350 131.440 67.670 131.760 ;
        RECT 67.750 131.440 68.070 131.760 ;
        RECT 68.150 131.440 68.470 131.760 ;
        RECT 89.145 131.440 89.465 131.760 ;
        RECT 89.545 131.440 89.865 131.760 ;
        RECT 89.945 131.440 90.265 131.760 ;
        RECT 90.345 131.440 90.665 131.760 ;
        RECT 111.340 131.440 111.660 131.760 ;
        RECT 111.740 131.440 112.060 131.760 ;
        RECT 112.140 131.440 112.460 131.760 ;
        RECT 112.540 131.440 112.860 131.760 ;
        RECT 133.535 131.440 133.855 131.760 ;
        RECT 133.935 131.440 134.255 131.760 ;
        RECT 134.335 131.440 134.655 131.760 ;
        RECT 134.735 131.440 135.055 131.760 ;
        RECT 66.950 126.000 67.270 126.320 ;
        RECT 67.350 126.000 67.670 126.320 ;
        RECT 67.750 126.000 68.070 126.320 ;
        RECT 68.150 126.000 68.470 126.320 ;
        RECT 89.145 126.000 89.465 126.320 ;
        RECT 89.545 126.000 89.865 126.320 ;
        RECT 89.945 126.000 90.265 126.320 ;
        RECT 90.345 126.000 90.665 126.320 ;
        RECT 111.340 126.000 111.660 126.320 ;
        RECT 111.740 126.000 112.060 126.320 ;
        RECT 112.140 126.000 112.460 126.320 ;
        RECT 112.540 126.000 112.860 126.320 ;
        RECT 133.535 126.000 133.855 126.320 ;
        RECT 133.935 126.000 134.255 126.320 ;
        RECT 134.335 126.000 134.655 126.320 ;
        RECT 134.735 126.000 135.055 126.320 ;
        RECT 66.950 120.560 67.270 120.880 ;
        RECT 67.350 120.560 67.670 120.880 ;
        RECT 67.750 120.560 68.070 120.880 ;
        RECT 68.150 120.560 68.470 120.880 ;
        RECT 89.145 120.560 89.465 120.880 ;
        RECT 89.545 120.560 89.865 120.880 ;
        RECT 89.945 120.560 90.265 120.880 ;
        RECT 90.345 120.560 90.665 120.880 ;
        RECT 111.340 120.560 111.660 120.880 ;
        RECT 111.740 120.560 112.060 120.880 ;
        RECT 112.140 120.560 112.460 120.880 ;
        RECT 112.540 120.560 112.860 120.880 ;
        RECT 133.535 120.560 133.855 120.880 ;
        RECT 133.935 120.560 134.255 120.880 ;
        RECT 134.335 120.560 134.655 120.880 ;
        RECT 134.735 120.560 135.055 120.880 ;
        RECT 66.950 115.120 67.270 115.440 ;
        RECT 67.350 115.120 67.670 115.440 ;
        RECT 67.750 115.120 68.070 115.440 ;
        RECT 68.150 115.120 68.470 115.440 ;
        RECT 89.145 115.120 89.465 115.440 ;
        RECT 89.545 115.120 89.865 115.440 ;
        RECT 89.945 115.120 90.265 115.440 ;
        RECT 90.345 115.120 90.665 115.440 ;
        RECT 111.340 115.120 111.660 115.440 ;
        RECT 111.740 115.120 112.060 115.440 ;
        RECT 112.140 115.120 112.460 115.440 ;
        RECT 112.540 115.120 112.860 115.440 ;
        RECT 133.535 115.120 133.855 115.440 ;
        RECT 133.935 115.120 134.255 115.440 ;
        RECT 134.335 115.120 134.655 115.440 ;
        RECT 134.735 115.120 135.055 115.440 ;
        RECT 66.950 109.680 67.270 110.000 ;
        RECT 67.350 109.680 67.670 110.000 ;
        RECT 67.750 109.680 68.070 110.000 ;
        RECT 68.150 109.680 68.470 110.000 ;
        RECT 89.145 109.680 89.465 110.000 ;
        RECT 89.545 109.680 89.865 110.000 ;
        RECT 89.945 109.680 90.265 110.000 ;
        RECT 90.345 109.680 90.665 110.000 ;
        RECT 111.340 109.680 111.660 110.000 ;
        RECT 111.740 109.680 112.060 110.000 ;
        RECT 112.140 109.680 112.460 110.000 ;
        RECT 112.540 109.680 112.860 110.000 ;
        RECT 133.535 109.680 133.855 110.000 ;
        RECT 133.935 109.680 134.255 110.000 ;
        RECT 134.335 109.680 134.655 110.000 ;
        RECT 134.735 109.680 135.055 110.000 ;
        RECT 66.950 104.240 67.270 104.560 ;
        RECT 67.350 104.240 67.670 104.560 ;
        RECT 67.750 104.240 68.070 104.560 ;
        RECT 68.150 104.240 68.470 104.560 ;
        RECT 89.145 104.240 89.465 104.560 ;
        RECT 89.545 104.240 89.865 104.560 ;
        RECT 89.945 104.240 90.265 104.560 ;
        RECT 90.345 104.240 90.665 104.560 ;
        RECT 111.340 104.240 111.660 104.560 ;
        RECT 111.740 104.240 112.060 104.560 ;
        RECT 112.140 104.240 112.460 104.560 ;
        RECT 112.540 104.240 112.860 104.560 ;
        RECT 133.535 104.240 133.855 104.560 ;
        RECT 133.935 104.240 134.255 104.560 ;
        RECT 134.335 104.240 134.655 104.560 ;
        RECT 134.735 104.240 135.055 104.560 ;
        RECT 66.950 98.800 67.270 99.120 ;
        RECT 67.350 98.800 67.670 99.120 ;
        RECT 67.750 98.800 68.070 99.120 ;
        RECT 68.150 98.800 68.470 99.120 ;
        RECT 89.145 98.800 89.465 99.120 ;
        RECT 89.545 98.800 89.865 99.120 ;
        RECT 89.945 98.800 90.265 99.120 ;
        RECT 90.345 98.800 90.665 99.120 ;
        RECT 111.340 98.800 111.660 99.120 ;
        RECT 111.740 98.800 112.060 99.120 ;
        RECT 112.140 98.800 112.460 99.120 ;
        RECT 112.540 98.800 112.860 99.120 ;
        RECT 133.535 98.800 133.855 99.120 ;
        RECT 133.935 98.800 134.255 99.120 ;
        RECT 134.335 98.800 134.655 99.120 ;
        RECT 134.735 98.800 135.055 99.120 ;
        RECT 66.950 93.360 67.270 93.680 ;
        RECT 67.350 93.360 67.670 93.680 ;
        RECT 67.750 93.360 68.070 93.680 ;
        RECT 68.150 93.360 68.470 93.680 ;
        RECT 89.145 93.360 89.465 93.680 ;
        RECT 89.545 93.360 89.865 93.680 ;
        RECT 89.945 93.360 90.265 93.680 ;
        RECT 90.345 93.360 90.665 93.680 ;
        RECT 111.340 93.360 111.660 93.680 ;
        RECT 111.740 93.360 112.060 93.680 ;
        RECT 112.140 93.360 112.460 93.680 ;
        RECT 112.540 93.360 112.860 93.680 ;
        RECT 133.535 93.360 133.855 93.680 ;
        RECT 133.935 93.360 134.255 93.680 ;
        RECT 134.335 93.360 134.655 93.680 ;
        RECT 134.735 93.360 135.055 93.680 ;
        RECT 66.950 87.920 67.270 88.240 ;
        RECT 67.350 87.920 67.670 88.240 ;
        RECT 67.750 87.920 68.070 88.240 ;
        RECT 68.150 87.920 68.470 88.240 ;
        RECT 89.145 87.920 89.465 88.240 ;
        RECT 89.545 87.920 89.865 88.240 ;
        RECT 89.945 87.920 90.265 88.240 ;
        RECT 90.345 87.920 90.665 88.240 ;
        RECT 111.340 87.920 111.660 88.240 ;
        RECT 111.740 87.920 112.060 88.240 ;
        RECT 112.140 87.920 112.460 88.240 ;
        RECT 112.540 87.920 112.860 88.240 ;
        RECT 133.535 87.920 133.855 88.240 ;
        RECT 133.935 87.920 134.255 88.240 ;
        RECT 134.335 87.920 134.655 88.240 ;
        RECT 134.735 87.920 135.055 88.240 ;
        RECT 66.950 82.480 67.270 82.800 ;
        RECT 67.350 82.480 67.670 82.800 ;
        RECT 67.750 82.480 68.070 82.800 ;
        RECT 68.150 82.480 68.470 82.800 ;
        RECT 89.145 82.480 89.465 82.800 ;
        RECT 89.545 82.480 89.865 82.800 ;
        RECT 89.945 82.480 90.265 82.800 ;
        RECT 90.345 82.480 90.665 82.800 ;
        RECT 111.340 82.480 111.660 82.800 ;
        RECT 111.740 82.480 112.060 82.800 ;
        RECT 112.140 82.480 112.460 82.800 ;
        RECT 112.540 82.480 112.860 82.800 ;
        RECT 133.535 82.480 133.855 82.800 ;
        RECT 133.935 82.480 134.255 82.800 ;
        RECT 134.335 82.480 134.655 82.800 ;
        RECT 134.735 82.480 135.055 82.800 ;
        RECT 66.950 77.040 67.270 77.360 ;
        RECT 67.350 77.040 67.670 77.360 ;
        RECT 67.750 77.040 68.070 77.360 ;
        RECT 68.150 77.040 68.470 77.360 ;
        RECT 89.145 77.040 89.465 77.360 ;
        RECT 89.545 77.040 89.865 77.360 ;
        RECT 89.945 77.040 90.265 77.360 ;
        RECT 90.345 77.040 90.665 77.360 ;
        RECT 111.340 77.040 111.660 77.360 ;
        RECT 111.740 77.040 112.060 77.360 ;
        RECT 112.140 77.040 112.460 77.360 ;
        RECT 112.540 77.040 112.860 77.360 ;
        RECT 133.535 77.040 133.855 77.360 ;
        RECT 133.935 77.040 134.255 77.360 ;
        RECT 134.335 77.040 134.655 77.360 ;
        RECT 134.735 77.040 135.055 77.360 ;
        RECT 66.950 71.600 67.270 71.920 ;
        RECT 67.350 71.600 67.670 71.920 ;
        RECT 67.750 71.600 68.070 71.920 ;
        RECT 68.150 71.600 68.470 71.920 ;
        RECT 89.145 71.600 89.465 71.920 ;
        RECT 89.545 71.600 89.865 71.920 ;
        RECT 89.945 71.600 90.265 71.920 ;
        RECT 90.345 71.600 90.665 71.920 ;
        RECT 111.340 71.600 111.660 71.920 ;
        RECT 111.740 71.600 112.060 71.920 ;
        RECT 112.140 71.600 112.460 71.920 ;
        RECT 112.540 71.600 112.860 71.920 ;
        RECT 133.535 71.600 133.855 71.920 ;
        RECT 133.935 71.600 134.255 71.920 ;
        RECT 134.335 71.600 134.655 71.920 ;
        RECT 134.735 71.600 135.055 71.920 ;
        RECT 66.950 66.160 67.270 66.480 ;
        RECT 67.350 66.160 67.670 66.480 ;
        RECT 67.750 66.160 68.070 66.480 ;
        RECT 68.150 66.160 68.470 66.480 ;
        RECT 89.145 66.160 89.465 66.480 ;
        RECT 89.545 66.160 89.865 66.480 ;
        RECT 89.945 66.160 90.265 66.480 ;
        RECT 90.345 66.160 90.665 66.480 ;
        RECT 111.340 66.160 111.660 66.480 ;
        RECT 111.740 66.160 112.060 66.480 ;
        RECT 112.140 66.160 112.460 66.480 ;
        RECT 112.540 66.160 112.860 66.480 ;
        RECT 133.535 66.160 133.855 66.480 ;
        RECT 133.935 66.160 134.255 66.480 ;
        RECT 134.335 66.160 134.655 66.480 ;
        RECT 134.735 66.160 135.055 66.480 ;
        RECT 66.950 60.720 67.270 61.040 ;
        RECT 67.350 60.720 67.670 61.040 ;
        RECT 67.750 60.720 68.070 61.040 ;
        RECT 68.150 60.720 68.470 61.040 ;
        RECT 89.145 60.720 89.465 61.040 ;
        RECT 89.545 60.720 89.865 61.040 ;
        RECT 89.945 60.720 90.265 61.040 ;
        RECT 90.345 60.720 90.665 61.040 ;
        RECT 111.340 60.720 111.660 61.040 ;
        RECT 111.740 60.720 112.060 61.040 ;
        RECT 112.140 60.720 112.460 61.040 ;
        RECT 112.540 60.720 112.860 61.040 ;
        RECT 133.535 60.720 133.855 61.040 ;
        RECT 133.935 60.720 134.255 61.040 ;
        RECT 134.335 60.720 134.655 61.040 ;
        RECT 134.735 60.720 135.055 61.040 ;
      LAYER met4 ;
        RECT 66.910 60.640 68.510 137.280 ;
        RECT 89.105 60.640 90.705 137.280 ;
        RECT 111.300 60.640 112.900 137.280 ;
        RECT 133.495 60.640 135.095 137.280 ;
    END
    PORT
      LAYER li1 ;
        RECT 47.005 103.045 47.345 103.415 ;
        RECT 47.005 99.945 47.345 100.315 ;
      LAYER mcon ;
        RECT 47.045 103.125 47.215 103.295 ;
        RECT 47.045 100.065 47.215 100.235 ;
      LAYER met1 ;
        RECT 43.750 103.280 44.070 103.340 ;
        RECT 46.985 103.280 47.275 103.325 ;
        RECT 43.750 103.140 47.275 103.280 ;
        RECT 43.750 103.080 44.070 103.140 ;
        RECT 46.985 103.095 47.275 103.140 ;
        RECT 46.985 100.220 47.275 100.265 ;
        RECT 53.870 100.220 54.190 100.280 ;
        RECT 46.985 100.080 54.190 100.220 ;
        RECT 46.985 100.035 47.275 100.080 ;
        RECT 53.870 100.020 54.190 100.080 ;
      LAYER via ;
        RECT 43.780 103.080 44.040 103.340 ;
        RECT 53.900 100.020 54.160 100.280 ;
      LAYER met2 ;
        RECT 43.780 103.050 44.040 103.370 ;
        RECT 43.840 101.525 43.980 103.050 ;
        RECT 43.770 101.155 44.050 101.525 ;
        RECT 53.900 99.990 54.160 100.310 ;
        RECT 53.960 98.125 54.100 99.990 ;
        RECT 53.890 97.755 54.170 98.125 ;
      LAYER via2 ;
        RECT 43.770 101.200 44.050 101.480 ;
        RECT 53.890 97.800 54.170 98.080 ;
      LAYER met3 ;
        RECT 28.510 101.640 29.470 101.790 ;
        RECT 28.510 101.490 42.000 101.640 ;
        RECT 43.745 101.490 44.075 101.505 ;
        RECT 28.510 101.190 44.075 101.490 ;
        RECT 28.510 101.040 42.000 101.190 ;
        RECT 43.745 101.175 44.075 101.190 ;
        RECT 28.510 100.890 29.470 101.040 ;
        RECT 34.530 98.240 35.490 98.390 ;
        RECT 34.530 98.090 42.000 98.240 ;
        RECT 53.865 98.090 54.195 98.105 ;
        RECT 34.530 97.790 54.195 98.090 ;
        RECT 34.530 97.640 42.000 97.790 ;
        RECT 53.865 97.775 54.195 97.790 ;
        RECT 34.530 97.490 35.490 97.640 ;
      LAYER via3 ;
        RECT 28.630 100.980 29.350 101.700 ;
        RECT 34.650 97.580 35.370 98.300 ;
      LAYER met4 ;
        RECT 4.000 220.470 6.000 220.760 ;
        RECT 30.670 220.470 30.970 225.760 ;
        RECT 33.430 220.470 33.730 225.760 ;
        RECT 36.190 220.470 36.490 225.760 ;
        RECT 38.950 220.470 39.250 225.760 ;
        RECT 41.710 220.470 42.010 225.760 ;
        RECT 44.470 220.470 44.770 225.760 ;
        RECT 47.230 220.470 47.530 225.760 ;
        RECT 49.990 220.470 50.290 225.760 ;
        RECT 52.750 220.470 53.050 225.760 ;
        RECT 55.510 220.470 55.810 225.760 ;
        RECT 58.270 220.470 58.570 225.760 ;
        RECT 61.030 220.470 61.330 225.760 ;
        RECT 63.790 220.470 64.090 225.760 ;
        RECT 66.550 220.470 66.850 225.760 ;
        RECT 69.310 220.470 69.610 225.760 ;
        RECT 72.070 220.470 72.370 225.760 ;
        RECT 4.000 218.470 81.820 220.470 ;
        RECT 4.000 56.210 6.000 218.470 ;
        RECT 28.535 101.790 29.445 101.795 ;
        RECT 23.700 100.890 33.660 101.790 ;
        RECT 23.700 56.210 24.600 100.890 ;
        RECT 28.535 100.885 29.445 100.890 ;
        RECT 34.555 98.370 35.465 98.395 ;
        RECT 32.690 97.470 37.110 98.370 ;
        RECT 32.690 56.210 33.590 97.470 ;
        RECT 4.000 54.210 100.360 56.210 ;
        RECT 4.000 5.000 6.000 54.210 ;
        RECT 23.700 42.880 24.600 54.210 ;
        RECT 32.690 51.260 33.590 54.210 ;
        RECT 32.690 50.360 133.390 51.260 ;
        RECT 23.700 41.980 114.070 42.880 ;
        RECT 113.170 0.000 114.070 41.980 ;
        RECT 132.490 0.000 133.390 50.360 ;
    END
  END VGND
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 45.665 136.955 45.835 137.125 ;
        RECT 47.045 136.955 47.215 137.125 ;
        RECT 52.565 136.955 52.735 137.125 ;
        RECT 58.080 136.985 58.200 137.095 ;
        RECT 59.005 136.955 59.175 137.125 ;
        RECT 64.525 136.955 64.695 137.125 ;
        RECT 70.045 136.955 70.215 137.125 ;
        RECT 71.885 136.955 72.055 137.125 ;
        RECT 77.405 136.955 77.575 137.125 ;
        RECT 82.925 136.955 83.095 137.125 ;
        RECT 84.765 136.955 84.935 137.125 ;
        RECT 90.285 136.955 90.455 137.125 ;
        RECT 95.805 136.955 95.975 137.125 ;
        RECT 97.645 136.955 97.815 137.125 ;
        RECT 103.165 136.955 103.335 137.125 ;
        RECT 108.685 136.955 108.855 137.125 ;
        RECT 110.525 136.955 110.695 137.125 ;
        RECT 116.045 136.955 116.215 137.125 ;
        RECT 121.565 136.955 121.735 137.125 ;
        RECT 123.405 136.955 123.575 137.125 ;
        RECT 128.925 136.955 129.095 137.125 ;
        RECT 132.600 136.985 132.720 137.095 ;
        RECT 133.985 136.955 134.155 137.125 ;
        RECT 45.665 131.515 45.835 131.685 ;
        RECT 47.045 131.515 47.215 131.685 ;
        RECT 52.565 131.515 52.735 131.685 ;
        RECT 58.085 131.655 58.255 131.685 ;
        RECT 58.080 131.545 58.255 131.655 ;
        RECT 58.085 131.515 58.255 131.545 ;
        RECT 59.005 131.515 59.175 131.685 ;
        RECT 63.605 131.515 63.775 131.685 ;
        RECT 64.525 131.515 64.695 131.685 ;
        RECT 69.125 131.515 69.295 131.685 ;
        RECT 70.045 131.515 70.215 131.685 ;
        RECT 70.960 131.545 71.080 131.655 ;
        RECT 71.885 131.515 72.055 131.685 ;
        RECT 75.565 131.515 75.735 131.685 ;
        RECT 77.405 131.515 77.575 131.685 ;
        RECT 81.085 131.515 81.255 131.685 ;
        RECT 82.925 131.515 83.095 131.685 ;
        RECT 83.840 131.545 83.960 131.655 ;
        RECT 84.765 131.515 84.935 131.685 ;
        RECT 88.445 131.515 88.615 131.685 ;
        RECT 90.285 131.515 90.455 131.685 ;
        RECT 93.965 131.515 94.135 131.685 ;
        RECT 95.805 131.515 95.975 131.685 ;
        RECT 96.720 131.545 96.840 131.655 ;
        RECT 97.645 131.515 97.815 131.685 ;
        RECT 101.325 131.515 101.495 131.685 ;
        RECT 103.165 131.515 103.335 131.685 ;
        RECT 106.845 131.515 107.015 131.685 ;
        RECT 108.685 131.515 108.855 131.685 ;
        RECT 109.600 131.545 109.720 131.655 ;
        RECT 110.525 131.515 110.695 131.685 ;
        RECT 114.205 131.515 114.375 131.685 ;
        RECT 116.045 131.515 116.215 131.685 ;
        RECT 119.725 131.515 119.895 131.685 ;
        RECT 121.565 131.515 121.735 131.685 ;
        RECT 122.480 131.545 122.600 131.655 ;
        RECT 123.405 131.515 123.575 131.685 ;
        RECT 127.085 131.515 127.255 131.685 ;
        RECT 128.925 131.515 129.095 131.685 ;
        RECT 132.600 131.545 132.720 131.655 ;
        RECT 133.985 131.515 134.155 131.685 ;
        RECT 45.665 126.075 45.835 126.245 ;
        RECT 47.045 126.075 47.215 126.245 ;
        RECT 52.565 126.075 52.735 126.245 ;
        RECT 58.085 126.215 58.255 126.245 ;
        RECT 58.080 126.105 58.255 126.215 ;
        RECT 58.085 126.075 58.255 126.105 ;
        RECT 59.005 126.075 59.175 126.245 ;
        RECT 63.605 126.075 63.775 126.245 ;
        RECT 64.525 126.075 64.695 126.245 ;
        RECT 69.125 126.075 69.295 126.245 ;
        RECT 70.045 126.075 70.215 126.245 ;
        RECT 70.960 126.105 71.080 126.215 ;
        RECT 71.885 126.075 72.055 126.245 ;
        RECT 75.565 126.075 75.735 126.245 ;
        RECT 77.405 126.075 77.575 126.245 ;
        RECT 81.085 126.075 81.255 126.245 ;
        RECT 82.925 126.075 83.095 126.245 ;
        RECT 83.840 126.105 83.960 126.215 ;
        RECT 84.765 126.075 84.935 126.245 ;
        RECT 88.445 126.075 88.615 126.245 ;
        RECT 90.285 126.075 90.455 126.245 ;
        RECT 93.965 126.075 94.135 126.245 ;
        RECT 95.805 126.075 95.975 126.245 ;
        RECT 96.720 126.105 96.840 126.215 ;
        RECT 97.645 126.075 97.815 126.245 ;
        RECT 101.325 126.075 101.495 126.245 ;
        RECT 103.165 126.075 103.335 126.245 ;
        RECT 106.845 126.075 107.015 126.245 ;
        RECT 108.685 126.075 108.855 126.245 ;
        RECT 109.600 126.105 109.720 126.215 ;
        RECT 110.525 126.075 110.695 126.245 ;
        RECT 114.205 126.075 114.375 126.245 ;
        RECT 116.045 126.075 116.215 126.245 ;
        RECT 119.725 126.075 119.895 126.245 ;
        RECT 121.565 126.075 121.735 126.245 ;
        RECT 122.480 126.105 122.600 126.215 ;
        RECT 123.405 126.075 123.575 126.245 ;
        RECT 127.085 126.075 127.255 126.245 ;
        RECT 128.925 126.075 129.095 126.245 ;
        RECT 132.600 126.105 132.720 126.215 ;
        RECT 133.985 126.075 134.155 126.245 ;
        RECT 45.665 120.635 45.835 120.805 ;
        RECT 47.045 120.635 47.215 120.805 ;
        RECT 52.565 120.635 52.735 120.805 ;
        RECT 58.085 120.775 58.255 120.805 ;
        RECT 58.080 120.665 58.255 120.775 ;
        RECT 58.085 120.635 58.255 120.665 ;
        RECT 59.005 120.635 59.175 120.805 ;
        RECT 63.605 120.635 63.775 120.805 ;
        RECT 64.525 120.635 64.695 120.805 ;
        RECT 69.125 120.635 69.295 120.805 ;
        RECT 70.045 120.635 70.215 120.805 ;
        RECT 70.960 120.665 71.080 120.775 ;
        RECT 71.885 120.635 72.055 120.805 ;
        RECT 75.565 120.635 75.735 120.805 ;
        RECT 77.405 120.635 77.575 120.805 ;
        RECT 81.085 120.635 81.255 120.805 ;
        RECT 82.925 120.635 83.095 120.805 ;
        RECT 83.840 120.665 83.960 120.775 ;
        RECT 84.765 120.635 84.935 120.805 ;
        RECT 88.445 120.635 88.615 120.805 ;
        RECT 90.285 120.635 90.455 120.805 ;
        RECT 93.965 120.635 94.135 120.805 ;
        RECT 95.805 120.635 95.975 120.805 ;
        RECT 96.720 120.665 96.840 120.775 ;
        RECT 97.645 120.635 97.815 120.805 ;
        RECT 101.325 120.635 101.495 120.805 ;
        RECT 103.165 120.635 103.335 120.805 ;
        RECT 106.845 120.635 107.015 120.805 ;
        RECT 108.685 120.635 108.855 120.805 ;
        RECT 109.600 120.665 109.720 120.775 ;
        RECT 110.525 120.635 110.695 120.805 ;
        RECT 114.205 120.635 114.375 120.805 ;
        RECT 116.045 120.635 116.215 120.805 ;
        RECT 119.725 120.635 119.895 120.805 ;
        RECT 121.565 120.635 121.735 120.805 ;
        RECT 122.480 120.665 122.600 120.775 ;
        RECT 123.405 120.635 123.575 120.805 ;
        RECT 127.085 120.635 127.255 120.805 ;
        RECT 128.925 120.635 129.095 120.805 ;
        RECT 132.600 120.665 132.720 120.775 ;
        RECT 133.985 120.635 134.155 120.805 ;
        RECT 45.665 115.195 45.835 115.365 ;
        RECT 47.045 115.195 47.215 115.365 ;
        RECT 52.565 115.195 52.735 115.365 ;
        RECT 58.085 115.335 58.255 115.365 ;
        RECT 58.080 115.225 58.255 115.335 ;
        RECT 58.085 115.195 58.255 115.225 ;
        RECT 59.005 115.195 59.175 115.365 ;
        RECT 63.605 115.195 63.775 115.365 ;
        RECT 64.525 115.195 64.695 115.365 ;
        RECT 69.125 115.195 69.295 115.365 ;
        RECT 70.045 115.195 70.215 115.365 ;
        RECT 70.960 115.225 71.080 115.335 ;
        RECT 71.885 115.195 72.055 115.365 ;
        RECT 75.565 115.195 75.735 115.365 ;
        RECT 77.405 115.195 77.575 115.365 ;
        RECT 81.085 115.195 81.255 115.365 ;
        RECT 82.925 115.195 83.095 115.365 ;
        RECT 83.840 115.225 83.960 115.335 ;
        RECT 84.765 115.195 84.935 115.365 ;
        RECT 88.445 115.195 88.615 115.365 ;
        RECT 90.285 115.195 90.455 115.365 ;
        RECT 93.965 115.195 94.135 115.365 ;
        RECT 95.805 115.195 95.975 115.365 ;
        RECT 96.720 115.225 96.840 115.335 ;
        RECT 97.645 115.195 97.815 115.365 ;
        RECT 101.325 115.195 101.495 115.365 ;
        RECT 103.165 115.195 103.335 115.365 ;
        RECT 106.845 115.195 107.015 115.365 ;
        RECT 108.685 115.195 108.855 115.365 ;
        RECT 109.600 115.225 109.720 115.335 ;
        RECT 110.525 115.195 110.695 115.365 ;
        RECT 114.205 115.195 114.375 115.365 ;
        RECT 116.045 115.195 116.215 115.365 ;
        RECT 119.725 115.195 119.895 115.365 ;
        RECT 121.565 115.195 121.735 115.365 ;
        RECT 122.480 115.225 122.600 115.335 ;
        RECT 123.405 115.195 123.575 115.365 ;
        RECT 127.085 115.195 127.255 115.365 ;
        RECT 128.925 115.195 129.095 115.365 ;
        RECT 132.600 115.225 132.720 115.335 ;
        RECT 133.985 115.195 134.155 115.365 ;
        RECT 45.665 109.755 45.835 109.925 ;
        RECT 47.045 109.755 47.215 109.925 ;
        RECT 52.565 109.755 52.735 109.925 ;
        RECT 58.085 109.895 58.255 109.925 ;
        RECT 58.080 109.785 58.255 109.895 ;
        RECT 58.085 109.755 58.255 109.785 ;
        RECT 59.005 109.755 59.175 109.925 ;
        RECT 59.920 109.785 60.040 109.895 ;
        RECT 60.385 109.755 60.555 109.925 ;
        RECT 61.765 109.755 61.935 109.925 ;
        RECT 63.605 109.755 63.775 109.925 ;
        RECT 64.525 109.755 64.695 109.925 ;
        RECT 69.125 109.755 69.295 109.925 ;
        RECT 70.045 109.755 70.215 109.925 ;
        RECT 70.960 109.785 71.080 109.895 ;
        RECT 71.885 109.755 72.055 109.925 ;
        RECT 75.565 109.755 75.735 109.925 ;
        RECT 77.405 109.755 77.575 109.925 ;
        RECT 81.085 109.755 81.255 109.925 ;
        RECT 82.925 109.755 83.095 109.925 ;
        RECT 83.840 109.785 83.960 109.895 ;
        RECT 84.765 109.755 84.935 109.925 ;
        RECT 88.445 109.755 88.615 109.925 ;
        RECT 90.285 109.755 90.455 109.925 ;
        RECT 93.965 109.755 94.135 109.925 ;
        RECT 95.805 109.755 95.975 109.925 ;
        RECT 96.720 109.785 96.840 109.895 ;
        RECT 97.645 109.755 97.815 109.925 ;
        RECT 101.325 109.755 101.495 109.925 ;
        RECT 103.165 109.755 103.335 109.925 ;
        RECT 106.845 109.755 107.015 109.925 ;
        RECT 108.685 109.755 108.855 109.925 ;
        RECT 109.600 109.785 109.720 109.895 ;
        RECT 110.525 109.755 110.695 109.925 ;
        RECT 114.205 109.755 114.375 109.925 ;
        RECT 116.045 109.755 116.215 109.925 ;
        RECT 119.725 109.755 119.895 109.925 ;
        RECT 121.565 109.755 121.735 109.925 ;
        RECT 122.480 109.785 122.600 109.895 ;
        RECT 123.405 109.755 123.575 109.925 ;
        RECT 127.085 109.755 127.255 109.925 ;
        RECT 128.925 109.755 129.095 109.925 ;
        RECT 132.600 109.785 132.720 109.895 ;
        RECT 133.985 109.755 134.155 109.925 ;
        RECT 45.665 104.315 45.835 104.485 ;
        RECT 47.045 104.315 47.225 104.485 ;
        RECT 48.425 104.315 48.595 104.485 ;
        RECT 50.720 104.345 50.840 104.455 ;
        RECT 52.105 104.315 52.275 104.485 ;
        RECT 52.560 104.315 52.730 104.485 ;
        RECT 53.955 104.340 54.115 104.450 ;
        RECT 54.870 104.315 55.040 104.485 ;
        RECT 57.160 104.315 57.340 104.485 ;
        RECT 57.635 104.350 57.795 104.460 ;
        RECT 59.005 104.315 59.175 104.485 ;
        RECT 61.305 104.315 61.475 104.485 ;
        RECT 64.525 104.315 64.695 104.485 ;
        RECT 66.825 104.315 66.995 104.485 ;
        RECT 70.045 104.315 70.215 104.485 ;
        RECT 70.515 104.340 70.675 104.450 ;
        RECT 71.885 104.315 72.055 104.485 ;
        RECT 75.565 104.315 75.735 104.485 ;
        RECT 77.405 104.315 77.575 104.485 ;
        RECT 81.085 104.315 81.255 104.485 ;
        RECT 82.925 104.315 83.095 104.485 ;
        RECT 83.840 104.345 83.960 104.455 ;
        RECT 84.765 104.315 84.935 104.485 ;
        RECT 88.445 104.315 88.615 104.485 ;
        RECT 90.285 104.315 90.455 104.485 ;
        RECT 93.965 104.315 94.135 104.485 ;
        RECT 95.805 104.315 95.975 104.485 ;
        RECT 96.720 104.345 96.840 104.455 ;
        RECT 97.645 104.315 97.815 104.485 ;
        RECT 101.325 104.315 101.495 104.485 ;
        RECT 103.165 104.315 103.335 104.485 ;
        RECT 106.845 104.315 107.015 104.485 ;
        RECT 108.685 104.315 108.855 104.485 ;
        RECT 109.600 104.345 109.720 104.455 ;
        RECT 110.525 104.315 110.695 104.485 ;
        RECT 114.205 104.315 114.375 104.485 ;
        RECT 116.045 104.315 116.215 104.485 ;
        RECT 119.725 104.315 119.895 104.485 ;
        RECT 121.565 104.315 121.735 104.485 ;
        RECT 122.480 104.345 122.600 104.455 ;
        RECT 123.405 104.315 123.575 104.485 ;
        RECT 127.085 104.315 127.255 104.485 ;
        RECT 128.925 104.315 129.095 104.485 ;
        RECT 132.600 104.345 132.720 104.455 ;
        RECT 133.985 104.315 134.155 104.485 ;
        RECT 45.665 98.875 45.835 99.045 ;
        RECT 47.045 98.875 47.225 99.045 ;
        RECT 48.425 98.875 48.595 99.045 ;
        RECT 52.565 98.875 52.735 99.045 ;
        RECT 53.945 98.875 54.115 99.045 ;
        RECT 55.320 98.905 55.440 99.015 ;
        RECT 55.785 98.875 55.955 99.045 ;
        RECT 57.165 98.875 57.335 99.045 ;
        RECT 57.635 98.910 57.795 99.020 ;
        RECT 59.005 98.875 59.175 99.045 ;
        RECT 62.685 98.875 62.855 99.045 ;
        RECT 64.525 98.875 64.695 99.045 ;
        RECT 68.205 98.875 68.375 99.045 ;
        RECT 70.045 98.875 70.215 99.045 ;
        RECT 70.960 98.905 71.080 99.015 ;
        RECT 71.885 98.875 72.055 99.045 ;
        RECT 75.565 98.875 75.735 99.045 ;
        RECT 77.405 98.875 77.575 99.045 ;
        RECT 81.085 98.875 81.255 99.045 ;
        RECT 82.925 98.875 83.095 99.045 ;
        RECT 83.840 98.905 83.960 99.015 ;
        RECT 84.765 98.875 84.935 99.045 ;
        RECT 88.445 98.875 88.615 99.045 ;
        RECT 90.285 98.875 90.455 99.045 ;
        RECT 93.965 98.875 94.135 99.045 ;
        RECT 95.805 98.875 95.975 99.045 ;
        RECT 96.720 98.905 96.840 99.015 ;
        RECT 97.645 98.875 97.815 99.045 ;
        RECT 101.325 98.875 101.495 99.045 ;
        RECT 103.165 98.875 103.335 99.045 ;
        RECT 106.845 98.875 107.015 99.045 ;
        RECT 108.685 98.875 108.855 99.045 ;
        RECT 109.600 98.905 109.720 99.015 ;
        RECT 110.525 98.875 110.695 99.045 ;
        RECT 114.205 98.875 114.375 99.045 ;
        RECT 116.045 98.875 116.215 99.045 ;
        RECT 119.725 98.875 119.895 99.045 ;
        RECT 121.565 98.875 121.735 99.045 ;
        RECT 122.480 98.905 122.600 99.015 ;
        RECT 123.405 98.875 123.575 99.045 ;
        RECT 127.085 98.875 127.255 99.045 ;
        RECT 128.925 98.875 129.095 99.045 ;
        RECT 132.600 98.905 132.720 99.015 ;
        RECT 133.985 98.875 134.155 99.045 ;
        RECT 45.665 93.435 45.835 93.605 ;
        RECT 47.045 93.435 47.215 93.605 ;
        RECT 50.735 93.460 50.895 93.570 ;
        RECT 52.565 93.435 52.735 93.605 ;
        RECT 55.050 93.435 55.220 93.605 ;
        RECT 56.060 93.435 56.230 93.605 ;
        RECT 56.240 93.465 56.360 93.575 ;
        RECT 57.630 93.435 57.800 93.605 ;
        RECT 58.080 93.465 58.200 93.575 ;
        RECT 59.005 93.435 59.175 93.605 ;
        RECT 59.925 93.435 60.095 93.605 ;
        RECT 61.305 93.435 61.475 93.605 ;
        RECT 62.685 93.435 62.855 93.605 ;
        RECT 64.525 93.435 64.695 93.605 ;
        RECT 68.205 93.435 68.375 93.605 ;
        RECT 70.045 93.435 70.215 93.605 ;
        RECT 70.960 93.465 71.080 93.575 ;
        RECT 71.885 93.435 72.055 93.605 ;
        RECT 75.565 93.435 75.735 93.605 ;
        RECT 77.405 93.435 77.575 93.605 ;
        RECT 81.085 93.435 81.255 93.605 ;
        RECT 82.925 93.435 83.095 93.605 ;
        RECT 83.840 93.465 83.960 93.575 ;
        RECT 84.765 93.435 84.935 93.605 ;
        RECT 88.445 93.435 88.615 93.605 ;
        RECT 90.285 93.435 90.455 93.605 ;
        RECT 93.965 93.435 94.135 93.605 ;
        RECT 95.805 93.435 95.975 93.605 ;
        RECT 96.720 93.465 96.840 93.575 ;
        RECT 97.645 93.435 97.815 93.605 ;
        RECT 101.325 93.435 101.495 93.605 ;
        RECT 103.165 93.435 103.335 93.605 ;
        RECT 106.845 93.435 107.015 93.605 ;
        RECT 108.685 93.435 108.855 93.605 ;
        RECT 109.600 93.465 109.720 93.575 ;
        RECT 110.525 93.435 110.695 93.605 ;
        RECT 114.205 93.435 114.375 93.605 ;
        RECT 116.045 93.435 116.215 93.605 ;
        RECT 119.725 93.435 119.895 93.605 ;
        RECT 121.565 93.435 121.735 93.605 ;
        RECT 122.480 93.465 122.600 93.575 ;
        RECT 123.405 93.435 123.575 93.605 ;
        RECT 127.085 93.435 127.255 93.605 ;
        RECT 128.925 93.435 129.095 93.605 ;
        RECT 132.600 93.465 132.720 93.575 ;
        RECT 133.985 93.435 134.155 93.605 ;
        RECT 45.665 87.995 45.835 88.165 ;
        RECT 47.045 87.995 47.215 88.165 ;
        RECT 52.565 87.995 52.735 88.165 ;
        RECT 55.335 87.995 55.505 88.165 ;
        RECT 56.705 87.995 56.875 88.165 ;
        RECT 58.085 88.135 58.255 88.165 ;
        RECT 58.080 88.025 58.255 88.135 ;
        RECT 58.085 87.995 58.255 88.025 ;
        RECT 59.005 87.995 59.175 88.165 ;
        RECT 63.605 87.995 63.775 88.165 ;
        RECT 64.525 87.995 64.695 88.165 ;
        RECT 69.125 87.995 69.295 88.165 ;
        RECT 70.045 87.995 70.215 88.165 ;
        RECT 70.960 88.025 71.080 88.135 ;
        RECT 71.885 87.995 72.055 88.165 ;
        RECT 75.565 87.995 75.735 88.165 ;
        RECT 77.405 87.995 77.575 88.165 ;
        RECT 81.085 87.995 81.255 88.165 ;
        RECT 82.925 87.995 83.095 88.165 ;
        RECT 83.840 88.025 83.960 88.135 ;
        RECT 84.765 87.995 84.935 88.165 ;
        RECT 88.445 87.995 88.615 88.165 ;
        RECT 90.285 87.995 90.455 88.165 ;
        RECT 93.965 87.995 94.135 88.165 ;
        RECT 95.805 87.995 95.975 88.165 ;
        RECT 96.720 88.025 96.840 88.135 ;
        RECT 97.645 87.995 97.815 88.165 ;
        RECT 101.325 87.995 101.495 88.165 ;
        RECT 103.165 87.995 103.335 88.165 ;
        RECT 106.845 87.995 107.015 88.165 ;
        RECT 108.685 87.995 108.855 88.165 ;
        RECT 109.600 88.025 109.720 88.135 ;
        RECT 110.525 87.995 110.695 88.165 ;
        RECT 114.205 87.995 114.375 88.165 ;
        RECT 116.045 87.995 116.215 88.165 ;
        RECT 119.725 87.995 119.895 88.165 ;
        RECT 121.565 87.995 121.735 88.165 ;
        RECT 122.480 88.025 122.600 88.135 ;
        RECT 123.405 87.995 123.575 88.165 ;
        RECT 127.085 87.995 127.255 88.165 ;
        RECT 128.925 87.995 129.095 88.165 ;
        RECT 132.600 88.025 132.720 88.135 ;
        RECT 133.985 87.995 134.155 88.165 ;
        RECT 45.665 82.555 45.835 82.725 ;
        RECT 47.045 82.555 47.215 82.725 ;
        RECT 52.565 82.555 52.735 82.725 ;
        RECT 58.085 82.695 58.255 82.725 ;
        RECT 58.080 82.585 58.255 82.695 ;
        RECT 58.085 82.555 58.255 82.585 ;
        RECT 59.005 82.555 59.175 82.725 ;
        RECT 63.605 82.555 63.775 82.725 ;
        RECT 64.525 82.555 64.695 82.725 ;
        RECT 69.125 82.555 69.295 82.725 ;
        RECT 70.045 82.555 70.215 82.725 ;
        RECT 70.960 82.585 71.080 82.695 ;
        RECT 71.885 82.555 72.055 82.725 ;
        RECT 75.565 82.555 75.735 82.725 ;
        RECT 77.405 82.555 77.575 82.725 ;
        RECT 81.085 82.555 81.255 82.725 ;
        RECT 82.925 82.555 83.095 82.725 ;
        RECT 83.840 82.585 83.960 82.695 ;
        RECT 84.765 82.555 84.935 82.725 ;
        RECT 88.445 82.555 88.615 82.725 ;
        RECT 90.285 82.555 90.455 82.725 ;
        RECT 93.965 82.555 94.135 82.725 ;
        RECT 95.805 82.555 95.975 82.725 ;
        RECT 96.720 82.585 96.840 82.695 ;
        RECT 97.645 82.555 97.815 82.725 ;
        RECT 101.325 82.555 101.495 82.725 ;
        RECT 103.165 82.555 103.335 82.725 ;
        RECT 106.845 82.555 107.015 82.725 ;
        RECT 108.685 82.555 108.855 82.725 ;
        RECT 109.600 82.585 109.720 82.695 ;
        RECT 110.525 82.555 110.695 82.725 ;
        RECT 114.205 82.555 114.375 82.725 ;
        RECT 116.045 82.555 116.215 82.725 ;
        RECT 119.725 82.555 119.895 82.725 ;
        RECT 121.565 82.555 121.735 82.725 ;
        RECT 122.480 82.585 122.600 82.695 ;
        RECT 123.405 82.555 123.575 82.725 ;
        RECT 127.085 82.555 127.255 82.725 ;
        RECT 128.925 82.555 129.095 82.725 ;
        RECT 132.600 82.585 132.720 82.695 ;
        RECT 133.985 82.555 134.155 82.725 ;
        RECT 45.665 77.115 45.835 77.285 ;
        RECT 47.045 77.115 47.215 77.285 ;
        RECT 52.565 77.115 52.735 77.285 ;
        RECT 58.085 77.255 58.255 77.285 ;
        RECT 58.080 77.145 58.255 77.255 ;
        RECT 58.085 77.115 58.255 77.145 ;
        RECT 59.005 77.115 59.175 77.285 ;
        RECT 63.605 77.115 63.775 77.285 ;
        RECT 64.525 77.115 64.695 77.285 ;
        RECT 69.125 77.115 69.295 77.285 ;
        RECT 70.045 77.115 70.215 77.285 ;
        RECT 70.960 77.145 71.080 77.255 ;
        RECT 71.885 77.115 72.055 77.285 ;
        RECT 75.565 77.115 75.735 77.285 ;
        RECT 77.405 77.115 77.575 77.285 ;
        RECT 81.085 77.115 81.255 77.285 ;
        RECT 82.925 77.115 83.095 77.285 ;
        RECT 83.840 77.145 83.960 77.255 ;
        RECT 84.765 77.115 84.935 77.285 ;
        RECT 88.445 77.115 88.615 77.285 ;
        RECT 90.285 77.115 90.455 77.285 ;
        RECT 93.965 77.115 94.135 77.285 ;
        RECT 95.805 77.115 95.975 77.285 ;
        RECT 96.720 77.145 96.840 77.255 ;
        RECT 97.645 77.115 97.815 77.285 ;
        RECT 101.325 77.115 101.495 77.285 ;
        RECT 103.165 77.115 103.335 77.285 ;
        RECT 106.845 77.115 107.015 77.285 ;
        RECT 108.685 77.115 108.855 77.285 ;
        RECT 109.600 77.145 109.720 77.255 ;
        RECT 110.525 77.115 110.695 77.285 ;
        RECT 114.205 77.115 114.375 77.285 ;
        RECT 116.045 77.115 116.215 77.285 ;
        RECT 119.725 77.115 119.895 77.285 ;
        RECT 121.565 77.115 121.735 77.285 ;
        RECT 122.480 77.145 122.600 77.255 ;
        RECT 123.405 77.115 123.575 77.285 ;
        RECT 127.085 77.115 127.255 77.285 ;
        RECT 128.925 77.115 129.095 77.285 ;
        RECT 132.600 77.145 132.720 77.255 ;
        RECT 133.985 77.115 134.155 77.285 ;
        RECT 45.665 71.675 45.835 71.845 ;
        RECT 47.045 71.675 47.215 71.845 ;
        RECT 52.565 71.675 52.735 71.845 ;
        RECT 58.085 71.815 58.255 71.845 ;
        RECT 58.080 71.705 58.255 71.815 ;
        RECT 58.085 71.675 58.255 71.705 ;
        RECT 59.005 71.675 59.175 71.845 ;
        RECT 63.605 71.675 63.775 71.845 ;
        RECT 64.525 71.675 64.695 71.845 ;
        RECT 69.125 71.675 69.295 71.845 ;
        RECT 70.045 71.675 70.215 71.845 ;
        RECT 70.960 71.705 71.080 71.815 ;
        RECT 71.885 71.675 72.055 71.845 ;
        RECT 75.565 71.675 75.735 71.845 ;
        RECT 77.405 71.675 77.575 71.845 ;
        RECT 81.085 71.675 81.255 71.845 ;
        RECT 82.925 71.675 83.095 71.845 ;
        RECT 83.840 71.705 83.960 71.815 ;
        RECT 84.765 71.675 84.935 71.845 ;
        RECT 88.445 71.675 88.615 71.845 ;
        RECT 90.285 71.675 90.455 71.845 ;
        RECT 93.965 71.675 94.135 71.845 ;
        RECT 95.805 71.675 95.975 71.845 ;
        RECT 96.720 71.705 96.840 71.815 ;
        RECT 97.645 71.675 97.815 71.845 ;
        RECT 101.325 71.675 101.495 71.845 ;
        RECT 103.165 71.675 103.335 71.845 ;
        RECT 106.845 71.675 107.015 71.845 ;
        RECT 108.685 71.675 108.855 71.845 ;
        RECT 109.600 71.705 109.720 71.815 ;
        RECT 110.525 71.675 110.695 71.845 ;
        RECT 114.205 71.675 114.375 71.845 ;
        RECT 116.045 71.675 116.215 71.845 ;
        RECT 119.725 71.675 119.895 71.845 ;
        RECT 121.565 71.675 121.735 71.845 ;
        RECT 122.480 71.705 122.600 71.815 ;
        RECT 123.405 71.675 123.575 71.845 ;
        RECT 127.085 71.675 127.255 71.845 ;
        RECT 128.925 71.675 129.095 71.845 ;
        RECT 132.600 71.705 132.720 71.815 ;
        RECT 133.985 71.675 134.155 71.845 ;
        RECT 45.665 66.235 45.835 66.405 ;
        RECT 47.045 66.235 47.215 66.405 ;
        RECT 52.565 66.235 52.735 66.405 ;
        RECT 58.085 66.375 58.255 66.405 ;
        RECT 58.080 66.265 58.255 66.375 ;
        RECT 58.085 66.235 58.255 66.265 ;
        RECT 59.005 66.235 59.175 66.405 ;
        RECT 63.605 66.235 63.775 66.405 ;
        RECT 64.525 66.235 64.695 66.405 ;
        RECT 69.125 66.235 69.295 66.405 ;
        RECT 70.045 66.235 70.215 66.405 ;
        RECT 70.960 66.265 71.080 66.375 ;
        RECT 71.885 66.235 72.055 66.405 ;
        RECT 75.565 66.235 75.735 66.405 ;
        RECT 77.405 66.235 77.575 66.405 ;
        RECT 81.085 66.235 81.255 66.405 ;
        RECT 82.925 66.235 83.095 66.405 ;
        RECT 83.840 66.265 83.960 66.375 ;
        RECT 84.765 66.235 84.935 66.405 ;
        RECT 88.445 66.235 88.615 66.405 ;
        RECT 90.285 66.235 90.455 66.405 ;
        RECT 93.965 66.235 94.135 66.405 ;
        RECT 95.805 66.235 95.975 66.405 ;
        RECT 96.720 66.265 96.840 66.375 ;
        RECT 97.645 66.235 97.815 66.405 ;
        RECT 101.325 66.235 101.495 66.405 ;
        RECT 103.165 66.235 103.335 66.405 ;
        RECT 106.845 66.235 107.015 66.405 ;
        RECT 108.685 66.235 108.855 66.405 ;
        RECT 109.600 66.265 109.720 66.375 ;
        RECT 110.525 66.235 110.695 66.405 ;
        RECT 114.205 66.235 114.375 66.405 ;
        RECT 116.045 66.235 116.215 66.405 ;
        RECT 119.725 66.235 119.895 66.405 ;
        RECT 121.565 66.235 121.735 66.405 ;
        RECT 122.480 66.265 122.600 66.375 ;
        RECT 123.405 66.235 123.575 66.405 ;
        RECT 127.085 66.235 127.255 66.405 ;
        RECT 128.925 66.235 129.095 66.405 ;
        RECT 132.600 66.265 132.720 66.375 ;
        RECT 133.985 66.235 134.155 66.405 ;
        RECT 45.665 60.795 45.835 60.965 ;
        RECT 47.045 60.795 47.215 60.965 ;
        RECT 52.565 60.795 52.735 60.965 ;
        RECT 58.080 60.825 58.200 60.935 ;
        RECT 59.005 60.795 59.175 60.965 ;
        RECT 64.525 60.795 64.695 60.965 ;
        RECT 70.045 60.795 70.215 60.965 ;
        RECT 71.885 60.795 72.055 60.965 ;
        RECT 77.405 60.795 77.575 60.965 ;
        RECT 82.925 60.795 83.095 60.965 ;
        RECT 84.765 60.795 84.935 60.965 ;
        RECT 90.285 60.795 90.455 60.965 ;
        RECT 95.805 60.795 95.975 60.965 ;
        RECT 97.645 60.795 97.815 60.965 ;
        RECT 103.165 60.795 103.335 60.965 ;
        RECT 108.685 60.795 108.855 60.965 ;
        RECT 110.525 60.795 110.695 60.965 ;
        RECT 116.045 60.795 116.215 60.965 ;
        RECT 121.565 60.795 121.735 60.965 ;
        RECT 123.405 60.795 123.575 60.965 ;
        RECT 128.925 60.795 129.095 60.965 ;
        RECT 132.600 60.825 132.720 60.935 ;
        RECT 133.985 60.795 134.155 60.965 ;
      LAYER li1 ;
        RECT 60.765 108.955 61.095 109.585 ;
        RECT 61.795 109.205 61.965 109.585 ;
        RECT 61.795 109.035 62.510 109.205 ;
        RECT 60.345 108.515 60.675 108.765 ;
        RECT 60.845 108.355 61.095 108.955 ;
        RECT 61.705 108.485 62.060 108.855 ;
        RECT 62.340 108.845 62.510 109.035 ;
        RECT 62.680 109.010 62.935 109.585 ;
        RECT 62.340 108.515 62.595 108.845 ;
        RECT 60.765 107.375 61.095 108.355 ;
        RECT 62.340 108.305 62.510 108.515 ;
        RECT 61.795 108.135 62.510 108.305 ;
        RECT 62.765 108.280 62.935 109.010 ;
        RECT 61.795 107.375 61.965 108.135 ;
        RECT 62.680 107.375 62.935 108.280 ;
        RECT 51.565 105.885 51.895 106.865 ;
        RECT 52.955 105.885 53.285 106.865 ;
        RECT 56.210 106.405 56.465 106.860 ;
        RECT 57.135 106.405 57.395 106.865 ;
        RECT 55.675 106.200 56.465 106.405 ;
        RECT 51.565 105.285 51.815 105.885 ;
        RECT 53.020 105.845 53.195 105.885 ;
        RECT 51.985 105.475 52.315 105.725 ;
        RECT 52.515 105.455 52.850 105.725 ;
        RECT 53.020 105.285 53.190 105.845 ;
        RECT 55.675 105.725 56.070 106.200 ;
        RECT 56.740 106.185 57.395 106.405 ;
        RECT 53.360 105.475 53.695 105.725 ;
        RECT 54.395 105.395 54.775 105.725 ;
        RECT 54.945 105.475 56.070 105.725 ;
        RECT 56.240 105.475 56.570 106.030 ;
        RECT 54.525 105.305 54.775 105.395 ;
        RECT 51.565 104.655 51.895 105.285 ;
        RECT 53.020 104.655 53.715 105.285 ;
        RECT 54.525 105.135 55.625 105.305 ;
        RECT 55.455 104.865 55.625 105.135 ;
        RECT 55.795 105.285 56.070 105.475 ;
        RECT 55.795 105.035 56.125 105.285 ;
        RECT 56.740 105.225 56.955 106.185 ;
        RECT 57.125 105.395 57.395 106.015 ;
        RECT 56.295 105.015 57.395 105.225 ;
        RECT 56.295 104.865 56.465 105.015 ;
        RECT 55.455 104.655 56.465 104.865 ;
        RECT 57.135 104.680 57.395 105.015 ;
        RECT 47.075 103.765 47.245 104.145 ;
        RECT 47.075 103.595 47.740 103.765 ;
        RECT 47.935 103.640 48.195 104.145 ;
        RECT 47.570 103.340 47.740 103.595 ;
        RECT 47.570 103.010 47.845 103.340 ;
        RECT 47.570 102.865 47.740 103.010 ;
        RECT 47.065 102.695 47.740 102.865 ;
        RECT 48.015 102.840 48.195 103.640 ;
        RECT 54.805 103.685 55.145 104.145 ;
        RECT 55.655 103.935 56.825 104.145 ;
        RECT 55.655 103.685 55.905 103.935 ;
        RECT 56.495 103.915 56.825 103.935 ;
        RECT 57.105 103.785 57.365 104.120 ;
        RECT 58.040 103.805 58.750 104.145 ;
        RECT 54.805 103.515 55.905 103.685 ;
        RECT 56.075 103.495 56.935 103.745 ;
        RECT 54.805 103.075 55.565 103.325 ;
        RECT 55.735 103.075 56.485 103.325 ;
        RECT 56.655 102.905 56.935 103.495 ;
        RECT 47.065 101.935 47.245 102.695 ;
        RECT 47.925 101.935 48.195 102.840 ;
        RECT 55.235 102.735 56.935 102.905 ;
        RECT 55.235 101.935 55.565 102.735 ;
        RECT 56.075 101.935 56.405 102.735 ;
        RECT 57.105 102.555 57.340 103.785 ;
        RECT 57.510 102.725 57.800 103.635 ;
        RECT 57.970 103.125 58.300 103.635 ;
        RECT 58.470 103.375 58.750 103.805 ;
        RECT 58.920 103.745 59.190 104.145 ;
        RECT 59.860 103.935 61.070 104.125 ;
        RECT 59.860 103.745 60.145 103.935 ;
        RECT 58.920 103.545 60.145 103.745 ;
        RECT 60.315 103.545 61.075 103.765 ;
        RECT 58.470 103.125 59.985 103.375 ;
        RECT 60.265 103.125 60.675 103.375 ;
        RECT 58.470 102.955 58.755 103.125 ;
        RECT 60.845 102.955 61.075 103.545 ;
        RECT 58.140 102.635 58.755 102.955 ;
        RECT 58.925 102.775 61.075 102.955 ;
        RECT 58.925 102.635 60.645 102.775 ;
        RECT 57.105 101.935 57.365 102.555 ;
        RECT 58.140 101.935 58.430 102.635 ;
        RECT 58.620 102.295 60.145 102.465 ;
        RECT 58.620 101.935 58.830 102.295 ;
        RECT 59.500 102.105 60.145 102.295 ;
        RECT 60.315 102.275 60.645 102.635 ;
        RECT 60.815 102.105 61.075 102.605 ;
        RECT 59.500 101.935 61.075 102.105 ;
        RECT 47.065 100.665 47.245 101.425 ;
        RECT 47.065 100.495 47.740 100.665 ;
        RECT 47.925 100.520 48.195 101.425 ;
        RECT 47.570 100.350 47.740 100.495 ;
        RECT 47.570 100.020 47.845 100.350 ;
        RECT 47.570 99.765 47.740 100.020 ;
        RECT 47.075 99.595 47.740 99.765 ;
        RECT 48.015 99.720 48.195 100.520 ;
        RECT 47.075 99.215 47.245 99.595 ;
        RECT 47.935 99.215 48.195 99.720 ;
        RECT 55.815 98.325 55.985 98.705 ;
        RECT 55.815 98.155 56.480 98.325 ;
        RECT 56.675 98.200 56.935 98.705 ;
        RECT 55.745 97.605 56.075 97.975 ;
        RECT 56.310 97.900 56.480 98.155 ;
        RECT 56.310 97.570 56.595 97.900 ;
        RECT 56.310 97.425 56.480 97.570 ;
        RECT 55.815 97.255 56.480 97.425 ;
        RECT 56.765 97.400 56.935 98.200 ;
        RECT 55.815 96.495 55.985 97.255 ;
        RECT 56.665 96.495 56.935 97.400 ;
        RECT 57.075 95.005 57.405 95.985 ;
        RECT 56.665 94.595 57.000 94.845 ;
        RECT 57.170 94.405 57.340 95.005 ;
        RECT 57.510 94.575 57.845 94.845 ;
        RECT 56.645 93.775 57.340 94.405 ;
        RECT 51.860 92.625 52.105 93.230 ;
        RECT 51.585 92.455 52.815 92.625 ;
        RECT 51.585 91.645 51.925 92.455 ;
        RECT 52.095 91.890 52.845 92.080 ;
        RECT 51.585 91.235 52.100 91.645 ;
        RECT 52.675 91.225 52.845 91.890 ;
        RECT 53.015 91.905 53.205 93.265 ;
        RECT 53.375 93.095 53.650 93.265 ;
        RECT 53.375 92.925 53.655 93.095 ;
        RECT 53.375 92.105 53.650 92.925 ;
        RECT 53.840 92.900 54.370 93.265 ;
        RECT 54.195 92.865 54.370 92.900 ;
        RECT 53.855 91.905 54.025 92.705 ;
        RECT 53.015 91.735 54.025 91.905 ;
        RECT 54.195 92.695 55.125 92.865 ;
        RECT 55.295 92.695 55.550 93.265 ;
        RECT 54.195 91.565 54.365 92.695 ;
        RECT 54.955 92.525 55.125 92.695 ;
        RECT 53.240 91.395 54.365 91.565 ;
        RECT 54.535 92.195 54.730 92.525 ;
        RECT 54.955 92.195 55.210 92.525 ;
        RECT 54.535 91.225 54.705 92.195 ;
        RECT 55.380 92.025 55.550 92.695 ;
        RECT 52.675 91.055 54.705 91.225 ;
        RECT 55.215 91.055 55.550 92.025 ;
        RECT 55.730 92.695 55.985 93.265 ;
        RECT 56.910 92.900 57.440 93.265 ;
        RECT 56.910 92.865 57.085 92.900 ;
        RECT 56.155 92.695 57.085 92.865 ;
        RECT 55.730 92.025 55.900 92.695 ;
        RECT 56.155 92.525 56.325 92.695 ;
        RECT 56.070 92.195 56.325 92.525 ;
        RECT 56.550 92.195 56.745 92.525 ;
        RECT 55.730 91.055 56.065 92.025 ;
        RECT 56.575 91.225 56.745 92.195 ;
        RECT 56.915 91.565 57.085 92.695 ;
        RECT 57.255 91.905 57.425 92.705 ;
        RECT 57.630 92.415 57.905 93.265 ;
        RECT 57.625 92.245 57.905 92.415 ;
        RECT 57.630 92.105 57.905 92.245 ;
        RECT 58.075 91.905 58.265 93.265 ;
        RECT 59.175 92.625 59.420 93.230 ;
        RECT 60.305 92.635 60.635 93.265 ;
        RECT 61.685 92.635 62.015 93.265 ;
        RECT 58.465 92.455 59.695 92.625 ;
        RECT 57.255 91.735 58.265 91.905 ;
        RECT 58.435 91.890 59.185 92.080 ;
        RECT 56.915 91.395 58.040 91.565 ;
        RECT 58.435 91.225 58.605 91.890 ;
        RECT 59.355 91.645 59.695 92.455 ;
        RECT 59.885 92.195 60.215 92.445 ;
        RECT 60.385 92.035 60.635 92.635 ;
        RECT 61.265 92.195 61.595 92.445 ;
        RECT 61.765 92.035 62.015 92.635 ;
        RECT 59.180 91.235 59.695 91.645 ;
        RECT 56.575 91.055 58.605 91.225 ;
        RECT 60.305 91.055 60.635 92.035 ;
        RECT 61.685 91.055 62.015 92.035 ;
        RECT 55.345 89.785 55.525 90.545 ;
        RECT 55.345 89.615 56.020 89.785 ;
        RECT 56.205 89.640 56.475 90.545 ;
        RECT 55.850 89.470 56.020 89.615 ;
        RECT 55.285 89.065 55.625 89.435 ;
        RECT 55.850 89.140 56.125 89.470 ;
        RECT 55.850 88.885 56.020 89.140 ;
        RECT 55.355 88.715 56.020 88.885 ;
        RECT 56.295 88.840 56.475 89.640 ;
        RECT 57.085 89.565 57.415 90.545 ;
        RECT 56.665 89.155 56.995 89.405 ;
        RECT 57.165 88.965 57.415 89.565 ;
        RECT 55.355 88.335 55.525 88.715 ;
        RECT 56.215 88.335 56.475 88.840 ;
        RECT 57.085 88.335 57.415 88.965 ;
      LAYER mcon ;
        RECT 60.385 108.565 60.555 108.735 ;
        RECT 60.845 108.565 61.015 108.735 ;
        RECT 61.765 108.565 61.935 108.735 ;
        RECT 53.025 105.845 53.195 106.015 ;
        RECT 52.105 105.505 52.275 105.675 ;
        RECT 52.565 105.505 52.735 105.675 ;
        RECT 53.485 105.505 53.655 105.675 ;
        RECT 56.245 105.845 56.415 106.015 ;
        RECT 57.165 105.505 57.335 105.675 ;
        RECT 47.965 103.805 48.135 103.975 ;
        RECT 56.705 103.465 56.875 103.635 ;
        RECT 54.865 103.125 55.035 103.295 ;
        RECT 56.245 103.125 56.415 103.295 ;
        RECT 57.170 103.125 57.340 103.295 ;
        RECT 58.085 103.465 58.255 103.635 ;
        RECT 60.400 103.125 60.570 103.295 ;
        RECT 57.625 102.785 57.795 102.955 ;
        RECT 59.005 102.785 59.175 102.955 ;
        RECT 47.965 99.385 48.135 99.555 ;
        RECT 56.705 98.365 56.875 98.535 ;
        RECT 55.785 97.685 55.955 97.855 ;
        RECT 56.705 94.625 56.875 94.795 ;
        RECT 57.625 94.625 57.795 94.795 ;
        RECT 56.705 93.945 56.875 94.115 ;
        RECT 53.025 92.925 53.195 93.095 ;
        RECT 52.565 91.905 52.735 92.075 ;
        RECT 53.485 92.925 53.655 93.095 ;
        RECT 55.325 91.225 55.495 91.395 ;
        RECT 55.785 92.925 55.955 93.095 ;
        RECT 58.085 92.585 58.255 92.755 ;
        RECT 58.545 91.905 58.715 92.075 ;
        RECT 59.925 92.245 60.095 92.415 ;
        RECT 61.765 92.585 61.935 92.755 ;
        RECT 61.305 92.245 61.475 92.415 ;
        RECT 55.325 89.185 55.495 89.355 ;
        RECT 57.165 90.205 57.335 90.375 ;
        RECT 56.705 89.185 56.875 89.355 ;
      LAYER met1 ;
        RECT 58.930 108.720 59.250 108.780 ;
        RECT 60.325 108.720 60.615 108.765 ;
        RECT 58.930 108.580 60.615 108.720 ;
        RECT 58.930 108.520 59.250 108.580 ;
        RECT 60.325 108.535 60.615 108.580 ;
        RECT 60.785 108.720 61.075 108.765 ;
        RECT 61.705 108.720 61.995 108.765 ;
        RECT 60.785 108.580 61.995 108.720 ;
        RECT 60.785 108.535 61.075 108.580 ;
        RECT 61.705 108.535 61.995 108.580 ;
        RECT 52.965 106.000 53.255 106.045 ;
        RECT 56.185 106.000 56.475 106.045 ;
        RECT 52.965 105.860 56.475 106.000 ;
        RECT 52.965 105.815 53.255 105.860 ;
        RECT 56.185 105.815 56.475 105.860 ;
        RECT 52.030 105.660 52.350 105.720 ;
        RECT 52.505 105.660 52.795 105.705 ;
        RECT 52.030 105.520 52.795 105.660 ;
        RECT 52.030 105.460 52.350 105.520 ;
        RECT 52.505 105.475 52.795 105.520 ;
        RECT 53.425 105.660 53.715 105.705 ;
        RECT 55.250 105.660 55.570 105.720 ;
        RECT 53.425 105.520 55.570 105.660 ;
        RECT 53.425 105.475 53.715 105.520 ;
        RECT 55.250 105.460 55.570 105.520 ;
        RECT 57.105 105.660 57.395 105.705 ;
        RECT 57.550 105.660 57.870 105.720 ;
        RECT 57.105 105.520 57.870 105.660 ;
        RECT 57.105 105.475 57.395 105.520 ;
        RECT 57.550 105.460 57.870 105.520 ;
        RECT 47.905 103.960 48.195 104.005 ;
        RECT 52.030 103.960 52.350 104.020 ;
        RECT 47.905 103.820 52.350 103.960 ;
        RECT 47.905 103.775 48.195 103.820 ;
        RECT 52.030 103.760 52.350 103.820 ;
        RECT 52.120 103.280 52.260 103.760 ;
        RECT 56.645 103.620 56.935 103.665 ;
        RECT 58.025 103.620 58.315 103.665 ;
        RECT 58.470 103.620 58.790 103.680 ;
        RECT 56.645 103.480 58.790 103.620 ;
        RECT 56.645 103.435 56.935 103.480 ;
        RECT 58.025 103.435 58.315 103.480 ;
        RECT 58.470 103.420 58.790 103.480 ;
        RECT 54.805 103.280 55.095 103.325 ;
        RECT 52.120 103.140 55.095 103.280 ;
        RECT 54.805 103.095 55.095 103.140 ;
        RECT 55.250 103.280 55.570 103.340 ;
        RECT 56.185 103.280 56.475 103.325 ;
        RECT 55.250 103.140 56.475 103.280 ;
        RECT 55.250 103.080 55.570 103.140 ;
        RECT 56.185 103.095 56.475 103.140 ;
        RECT 57.105 103.280 57.400 103.325 ;
        RECT 60.340 103.280 60.630 103.325 ;
        RECT 57.105 103.140 60.630 103.280 ;
        RECT 57.105 103.095 57.400 103.140 ;
        RECT 60.340 103.095 60.630 103.140 ;
        RECT 56.260 102.600 56.400 103.095 ;
        RECT 57.550 102.740 57.870 103.000 ;
        RECT 58.930 102.740 59.250 103.000 ;
        RECT 59.020 102.600 59.160 102.740 ;
        RECT 56.260 102.460 59.160 102.600 ;
        RECT 47.905 99.540 48.195 99.585 ;
        RECT 53.410 99.540 53.730 99.600 ;
        RECT 47.905 99.400 53.730 99.540 ;
        RECT 47.905 99.355 48.195 99.400 ;
        RECT 53.410 99.340 53.730 99.400 ;
        RECT 56.645 98.520 56.935 98.565 ;
        RECT 57.550 98.520 57.870 98.580 ;
        RECT 56.645 98.380 57.870 98.520 ;
        RECT 56.645 98.335 56.935 98.380 ;
        RECT 57.550 98.320 57.870 98.380 ;
        RECT 55.250 97.840 55.570 97.900 ;
        RECT 55.725 97.840 56.015 97.885 ;
        RECT 55.250 97.700 56.015 97.840 ;
        RECT 55.250 97.640 55.570 97.700 ;
        RECT 55.725 97.655 56.015 97.700 ;
        RECT 53.410 94.780 53.730 94.840 ;
        RECT 56.645 94.780 56.935 94.825 ;
        RECT 53.410 94.640 56.935 94.780 ;
        RECT 53.410 94.580 53.730 94.640 ;
        RECT 56.645 94.595 56.935 94.640 ;
        RECT 57.565 94.780 57.855 94.825 ;
        RECT 58.930 94.780 59.250 94.840 ;
        RECT 57.565 94.640 59.250 94.780 ;
        RECT 57.565 94.595 57.855 94.640 ;
        RECT 58.930 94.580 59.250 94.640 ;
        RECT 52.950 94.100 53.270 94.160 ;
        RECT 56.645 94.100 56.935 94.145 ;
        RECT 61.230 94.100 61.550 94.160 ;
        RECT 52.950 93.960 61.550 94.100 ;
        RECT 52.950 93.900 53.270 93.960 ;
        RECT 56.645 93.915 56.935 93.960 ;
        RECT 61.230 93.900 61.550 93.960 ;
        RECT 52.950 92.880 53.270 93.140 ;
        RECT 53.410 92.880 53.730 93.140 ;
        RECT 55.250 93.080 55.570 93.140 ;
        RECT 55.725 93.080 56.015 93.125 ;
        RECT 55.250 92.940 56.015 93.080 ;
        RECT 55.250 92.880 55.570 92.940 ;
        RECT 55.725 92.895 56.015 92.940 ;
        RECT 58.025 92.740 58.315 92.785 ;
        RECT 61.705 92.740 61.995 92.785 ;
        RECT 58.025 92.600 61.995 92.740 ;
        RECT 58.025 92.555 58.315 92.600 ;
        RECT 61.705 92.555 61.995 92.600 ;
        RECT 57.550 92.200 57.870 92.460 ;
        RECT 59.865 92.400 60.155 92.445 ;
        RECT 58.560 92.260 60.155 92.400 ;
        RECT 58.560 92.120 58.700 92.260 ;
        RECT 59.865 92.215 60.155 92.260 ;
        RECT 61.230 92.200 61.550 92.460 ;
        RECT 52.505 92.060 52.795 92.105 ;
        RECT 58.470 92.060 58.790 92.120 ;
        RECT 52.505 91.920 58.790 92.060 ;
        RECT 52.505 91.875 52.795 91.920 ;
        RECT 58.470 91.860 58.790 91.920 ;
        RECT 55.250 91.180 55.570 91.440 ;
        RECT 57.105 90.360 57.395 90.405 ;
        RECT 57.550 90.360 57.870 90.420 ;
        RECT 57.105 90.220 57.870 90.360 ;
        RECT 57.105 90.175 57.395 90.220 ;
        RECT 57.550 90.160 57.870 90.220 ;
        RECT 53.870 89.680 54.190 89.740 ;
        RECT 53.870 89.540 56.860 89.680 ;
        RECT 53.870 89.480 54.190 89.540 ;
        RECT 55.250 89.140 55.570 89.400 ;
        RECT 56.720 89.385 56.860 89.540 ;
        RECT 56.645 89.155 56.935 89.385 ;
      LAYER via ;
        RECT 58.960 108.520 59.220 108.780 ;
        RECT 52.060 105.460 52.320 105.720 ;
        RECT 55.280 105.460 55.540 105.720 ;
        RECT 57.580 105.460 57.840 105.720 ;
        RECT 52.060 103.760 52.320 104.020 ;
        RECT 58.500 103.420 58.760 103.680 ;
        RECT 55.280 103.080 55.540 103.340 ;
        RECT 57.580 102.740 57.840 103.000 ;
        RECT 58.960 102.740 59.220 103.000 ;
        RECT 53.440 99.340 53.700 99.600 ;
        RECT 57.580 98.320 57.840 98.580 ;
        RECT 55.280 97.640 55.540 97.900 ;
        RECT 53.440 94.580 53.700 94.840 ;
        RECT 58.960 94.580 59.220 94.840 ;
        RECT 52.980 93.900 53.240 94.160 ;
        RECT 61.260 93.900 61.520 94.160 ;
        RECT 52.980 92.880 53.240 93.140 ;
        RECT 53.440 92.880 53.700 93.140 ;
        RECT 55.280 92.880 55.540 93.140 ;
        RECT 57.580 92.200 57.840 92.460 ;
        RECT 61.260 92.200 61.520 92.460 ;
        RECT 58.500 91.860 58.760 92.120 ;
        RECT 55.280 91.180 55.540 91.440 ;
        RECT 57.580 90.160 57.840 90.420 ;
        RECT 53.900 89.480 54.160 89.740 ;
        RECT 55.280 89.140 55.540 89.400 ;
      LAYER met2 ;
        RECT 58.960 108.490 59.220 108.810 ;
        RECT 52.060 105.430 52.320 105.750 ;
        RECT 55.280 105.430 55.540 105.750 ;
        RECT 57.580 105.430 57.840 105.750 ;
        RECT 52.120 104.050 52.260 105.430 ;
        RECT 52.060 103.730 52.320 104.050 ;
        RECT 55.340 103.370 55.480 105.430 ;
        RECT 55.280 103.050 55.540 103.370 ;
        RECT 57.640 103.030 57.780 105.430 ;
        RECT 58.500 103.390 58.760 103.710 ;
        RECT 57.580 102.710 57.840 103.030 ;
        RECT 53.440 99.310 53.700 99.630 ;
        RECT 53.500 94.870 53.640 99.310 ;
        RECT 57.640 98.610 57.780 102.710 ;
        RECT 57.580 98.290 57.840 98.610 ;
        RECT 55.280 97.610 55.540 97.930 ;
        RECT 53.440 94.550 53.700 94.870 ;
        RECT 52.980 93.870 53.240 94.190 ;
        RECT 53.040 93.170 53.180 93.870 ;
        RECT 53.500 93.170 53.640 94.550 ;
        RECT 55.340 93.170 55.480 97.610 ;
        RECT 52.980 92.850 53.240 93.170 ;
        RECT 53.440 92.850 53.700 93.170 ;
        RECT 55.280 92.850 55.540 93.170 ;
        RECT 53.500 91.890 53.640 92.850 ;
        RECT 57.580 92.170 57.840 92.490 ;
        RECT 53.500 91.750 54.100 91.890 ;
        RECT 53.960 89.770 54.100 91.750 ;
        RECT 55.280 91.150 55.540 91.470 ;
        RECT 53.900 89.450 54.160 89.770 ;
        RECT 55.340 89.430 55.480 91.150 ;
        RECT 57.640 90.450 57.780 92.170 ;
        RECT 58.560 92.150 58.700 103.390 ;
        RECT 59.020 103.030 59.160 108.490 ;
        RECT 58.960 102.710 59.220 103.030 ;
        RECT 59.020 94.870 59.160 102.710 ;
        RECT 58.960 94.550 59.220 94.870 ;
        RECT 61.260 93.870 61.520 94.190 ;
        RECT 61.320 92.490 61.460 93.870 ;
        RECT 61.260 92.170 61.520 92.490 ;
        RECT 58.500 91.830 58.760 92.150 ;
        RECT 57.580 90.130 57.840 90.450 ;
        RECT 55.280 89.110 55.540 89.430 ;
  END
END tt_um_DIGI_OTA
END LIBRARY

