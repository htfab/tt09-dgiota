VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_template
  CLASS BLOCK ;
  FOREIGN tt_um_template ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 142.830 224.760 143.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 145.590 224.760 145.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 140.070 224.760 140.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 53.560 209.800 54.155 209.805 ;
        RECT 53.560 209.465 55.165 209.800 ;
        RECT 53.560 208.145 53.735 209.465 ;
        RECT 53.560 207.595 54.155 208.145 ;
      LAYER mcon ;
        RECT 54.910 209.545 55.080 209.715 ;
      LAYER met1 ;
        RECT 54.830 215.930 65.715 216.075 ;
        RECT 54.830 215.740 65.725 215.930 ;
        RECT 54.830 209.830 55.165 215.740 ;
        RECT 65.365 214.920 65.725 215.740 ;
        RECT 54.800 209.435 55.195 209.830 ;
        RECT 54.830 209.385 55.165 209.435 ;
        RECT 65.360 97.845 65.735 189.265 ;
        RECT 65.330 97.470 65.765 97.845 ;
      LAYER via ;
        RECT 65.415 215.020 65.675 215.280 ;
        RECT 65.360 188.860 65.735 189.235 ;
        RECT 65.360 97.470 65.735 97.845 ;
      LAYER met2 ;
        RECT 65.360 189.235 65.735 215.435 ;
        RECT 65.330 188.860 65.765 189.235 ;
        RECT 65.360 188.800 65.735 188.860 ;
        RECT 65.360 23.320 65.735 97.875 ;
        RECT 65.315 22.945 65.780 23.320 ;
      LAYER via2 ;
        RECT 65.360 22.945 65.735 23.320 ;
      LAYER met3 ;
        RECT 65.335 23.315 65.760 23.345 ;
        RECT 65.335 23.140 107.990 23.315 ;
        RECT 65.335 22.940 151.615 23.140 ;
        RECT 65.335 22.920 65.760 22.940 ;
        RECT 107.100 22.765 151.615 22.940 ;
        RECT 150.690 0.280 151.590 22.765 ;
      LAYER via3 ;
        RECT 151.020 0.460 151.340 0.780 ;
      LAYER met4 ;
        RECT 150.810 0.000 151.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 24.190 197.255 25.390 197.495 ;
      LAYER mcon ;
        RECT 24.280 197.310 24.450 197.480 ;
      LAYER met1 ;
        RECT 20.305 200.755 24.490 201.005 ;
        RECT 19.540 199.475 19.860 199.480 ;
        RECT 20.305 199.475 20.555 200.755 ;
        RECT 19.540 199.225 20.555 199.475 ;
        RECT 19.540 199.220 19.860 199.225 ;
        RECT 24.240 197.245 24.490 200.755 ;
        RECT 19.540 182.970 19.860 183.090 ;
        RECT 19.540 182.570 19.870 182.970 ;
        RECT 19.540 182.330 19.860 182.570 ;
        RECT 19.570 181.400 19.835 182.330 ;
        RECT 19.575 114.030 19.825 181.400 ;
        RECT 19.540 113.770 19.860 114.030 ;
        RECT 19.575 113.745 19.825 113.770 ;
      LAYER via ;
        RECT 19.570 199.220 19.830 199.480 ;
        RECT 19.550 182.600 19.870 182.940 ;
        RECT 19.570 113.770 19.830 114.030 ;
      LAYER met2 ;
        RECT 19.570 199.190 19.830 199.510 ;
        RECT 19.575 183.600 19.825 199.190 ;
        RECT 19.530 182.940 19.870 183.600 ;
        RECT 19.520 182.600 19.900 182.940 ;
        RECT 19.530 182.540 19.870 182.600 ;
        RECT 19.375 12.835 20.025 114.145 ;
      LAYER via2 ;
        RECT 19.420 12.900 19.980 13.460 ;
      LAYER met3 ;
        RECT 19.210 13.470 20.820 13.500 ;
        RECT 19.210 12.910 132.340 13.470 ;
        RECT 19.210 12.880 20.820 12.910 ;
        RECT 19.395 12.875 20.005 12.880 ;
        RECT 131.780 0.130 132.340 12.910 ;
      LAYER via3 ;
        RECT 131.905 0.205 132.225 0.525 ;
      LAYER met4 ;
        RECT 131.490 0.000 132.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 23.850 213.395 24.315 213.445 ;
        RECT 23.850 213.185 24.950 213.395 ;
        RECT 23.850 213.140 24.315 213.185 ;
        RECT 24.620 213.155 24.950 213.185 ;
      LAYER mcon ;
        RECT 23.905 213.235 24.075 213.405 ;
      LAYER met1 ;
        RECT 9.985 216.905 10.765 216.945 ;
        RECT 9.985 216.655 23.455 216.905 ;
        RECT 9.985 216.615 10.765 216.655 ;
        RECT 23.205 213.445 23.455 216.655 ;
        RECT 23.840 213.445 24.145 213.475 ;
        RECT 23.205 213.195 24.345 213.445 ;
        RECT 23.840 213.170 24.145 213.195 ;
        RECT 10.070 124.645 10.465 186.475 ;
      LAYER via ;
        RECT 10.120 216.650 10.380 216.910 ;
        RECT 10.095 186.040 10.410 186.360 ;
        RECT 10.095 124.720 10.410 125.035 ;
      LAYER met2 ;
        RECT 10.095 186.835 10.410 216.955 ;
        RECT 10.080 185.945 10.425 186.835 ;
        RECT 10.095 7.270 10.410 125.095 ;
        RECT 15.865 7.270 16.225 7.370 ;
        RECT 10.095 6.955 16.315 7.270 ;
        RECT 15.865 6.920 16.225 6.955 ;
      LAYER via2 ;
        RECT 15.905 7.015 16.185 7.295 ;
      LAYER met3 ;
        RECT 15.800 7.400 112.955 7.410 ;
        RECT 15.800 6.920 113.120 7.400 ;
        RECT 112.115 0.180 113.120 6.920 ;
      LAYER via3 ;
        RECT 112.435 0.540 112.755 0.860 ;
      LAYER met4 ;
        RECT 112.170 0.000 113.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 92.850 0.000 93.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 73.530 0.000 74.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 54.210 0.000 55.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 34.890 0.000 35.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 15.570 0.000 16.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 137.310 224.760 137.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 134.550 224.760 134.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 131.790 224.760 132.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 129.030 224.760 129.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 126.270 224.760 126.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 123.510 224.760 123.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 120.750 224.760 121.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 117.990 224.760 118.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 115.230 224.760 115.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 112.470 224.760 112.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 109.710 224.760 110.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 106.950 224.760 107.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 104.190 224.760 104.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 101.430 224.760 101.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 98.670 224.760 98.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 95.910 224.760 96.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 48.990 224.760 49.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 46.230 224.760 46.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 43.470 224.760 43.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 40.710 224.760 41.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 37.950 224.760 38.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 35.190 224.760 35.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 32.430 224.760 32.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 29.670 224.760 29.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 71.070 224.760 71.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 68.310 224.760 68.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 65.550 224.760 65.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 62.790 224.760 63.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 60.030 224.760 60.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 57.270 224.760 57.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 54.510 224.760 54.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 51.750 224.760 52.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 93.150 224.760 93.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 90.390 224.760 90.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 87.630 224.760 87.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 84.870 224.760 85.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 82.110 224.760 82.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 79.350 224.760 79.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 76.590 224.760 76.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 73.830 224.760 74.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 0.223500 ;
    ANTENNADIFFAREA 5.549500 ;
    PORT
      LAYER nwell ;
        RECT 29.910 216.000 32.750 216.010 ;
        RECT 22.250 214.990 23.090 215.000 ;
        RECT 22.250 213.395 25.870 214.990 ;
        RECT 29.910 214.405 33.125 216.000 ;
        RECT 32.285 214.395 33.125 214.405 ;
        RECT 22.900 213.385 25.870 213.395 ;
        RECT 22.900 209.095 26.010 210.700 ;
        RECT 40.150 208.695 45.340 210.300 ;
        RECT 51.750 208.645 56.140 210.250 ;
        RECT 32.900 205.380 33.740 205.400 ;
        RECT 23.270 205.330 26.130 205.350 ;
        RECT 22.960 203.745 26.130 205.330 ;
        RECT 30.260 203.795 33.740 205.380 ;
        RECT 30.260 203.775 33.200 203.795 ;
        RECT 22.960 203.725 23.800 203.745 ;
        RECT 54.460 199.600 57.200 199.610 ;
        RECT 23.290 197.485 26.310 199.090 ;
        RECT 54.460 198.005 57.840 199.600 ;
        RECT 57.000 197.995 57.840 198.005 ;
        RECT 48.530 192.100 49.370 192.120 ;
        RECT 45.300 190.515 49.370 192.100 ;
        RECT 45.300 190.495 49.030 190.515 ;
      LAYER li1 ;
        RECT 30.100 215.735 31.480 215.905 ;
        RECT 22.440 214.725 22.900 214.895 ;
        RECT 22.525 213.560 22.815 214.725 ;
        RECT 24.300 214.715 25.680 214.885 ;
        RECT 24.640 213.575 24.850 214.715 ;
        RECT 31.055 214.595 31.385 215.735 ;
        RECT 32.475 215.725 32.935 215.895 ;
        RECT 32.560 214.560 32.850 215.725 ;
        RECT 23.090 210.425 23.550 210.595 ;
        RECT 24.440 210.425 25.820 210.595 ;
        RECT 23.175 209.260 23.465 210.425 ;
        RECT 24.780 209.285 24.990 210.425 ;
        RECT 40.340 210.025 43.560 210.195 ;
        RECT 44.690 210.025 45.150 210.195 ;
        RECT 41.395 209.175 41.565 210.025 ;
        RECT 42.235 209.515 42.405 210.025 ;
        RECT 44.775 208.860 45.065 210.025 ;
        RECT 51.940 209.975 54.240 210.145 ;
        RECT 55.490 209.975 55.950 210.145 ;
        RECT 52.455 209.575 53.390 209.975 ;
        RECT 55.575 208.810 55.865 209.975 ;
        RECT 23.150 205.055 23.610 205.225 ;
        RECT 24.560 205.075 25.940 205.245 ;
        RECT 30.450 205.105 31.830 205.275 ;
        RECT 33.090 205.125 33.550 205.295 ;
        RECT 23.235 203.890 23.525 205.055 ;
        RECT 24.900 203.935 25.110 205.075 ;
        RECT 31.405 203.965 31.735 205.105 ;
        RECT 33.175 203.960 33.465 205.125 ;
        RECT 54.650 199.335 56.030 199.505 ;
        RECT 23.480 198.815 23.940 198.985 ;
        RECT 24.740 198.815 26.120 198.985 ;
        RECT 23.565 197.650 23.855 198.815 ;
        RECT 25.080 197.675 25.290 198.815 ;
        RECT 54.990 198.195 55.200 199.335 ;
        RECT 57.190 199.325 57.650 199.495 ;
        RECT 55.370 198.185 55.700 199.165 ;
        RECT 55.470 197.815 55.700 198.185 ;
        RECT 57.275 198.160 57.565 199.325 ;
        RECT 55.470 197.585 56.865 197.815 ;
        RECT 55.370 196.955 55.700 197.585 ;
        RECT 45.490 191.825 47.790 191.995 ;
        RECT 48.720 191.845 49.180 192.015 ;
        RECT 46.005 191.425 46.940 191.825 ;
        RECT 45.575 190.895 46.035 190.915 ;
        RECT 44.370 190.435 46.035 190.895 ;
        RECT 48.805 190.680 49.095 191.845 ;
        RECT 44.370 190.170 45.230 190.435 ;
        RECT 45.575 190.185 46.035 190.435 ;
      LAYER mcon ;
        RECT 30.245 215.735 30.415 215.905 ;
        RECT 30.705 215.735 30.875 215.905 ;
        RECT 31.165 215.735 31.335 215.905 ;
        RECT 22.585 214.725 22.755 214.895 ;
        RECT 24.445 214.715 24.615 214.885 ;
        RECT 24.905 214.715 25.075 214.885 ;
        RECT 25.365 214.715 25.535 214.885 ;
        RECT 32.620 215.725 32.790 215.895 ;
        RECT 23.235 210.425 23.405 210.595 ;
        RECT 24.585 210.425 24.755 210.595 ;
        RECT 25.045 210.425 25.215 210.595 ;
        RECT 25.505 210.425 25.675 210.595 ;
        RECT 40.485 210.025 40.655 210.195 ;
        RECT 40.945 210.025 41.115 210.195 ;
        RECT 41.405 210.025 41.575 210.195 ;
        RECT 41.865 210.025 42.035 210.195 ;
        RECT 42.325 210.025 42.495 210.195 ;
        RECT 42.785 210.025 42.955 210.195 ;
        RECT 43.245 210.025 43.415 210.195 ;
        RECT 44.835 210.025 45.005 210.195 ;
        RECT 52.085 209.975 52.255 210.145 ;
        RECT 52.545 209.975 52.715 210.145 ;
        RECT 53.005 209.975 53.175 210.145 ;
        RECT 53.465 209.975 53.635 210.145 ;
        RECT 53.925 209.975 54.095 210.145 ;
        RECT 55.635 209.975 55.805 210.145 ;
        RECT 23.295 205.055 23.465 205.225 ;
        RECT 24.705 205.075 24.875 205.245 ;
        RECT 25.165 205.075 25.335 205.245 ;
        RECT 25.625 205.075 25.795 205.245 ;
        RECT 30.595 205.105 30.765 205.275 ;
        RECT 31.055 205.105 31.225 205.275 ;
        RECT 31.515 205.105 31.685 205.275 ;
        RECT 33.235 205.125 33.405 205.295 ;
        RECT 54.795 199.335 54.965 199.505 ;
        RECT 55.255 199.335 55.425 199.505 ;
        RECT 55.715 199.335 55.885 199.505 ;
        RECT 23.625 198.815 23.795 198.985 ;
        RECT 24.885 198.815 25.055 198.985 ;
        RECT 25.345 198.815 25.515 198.985 ;
        RECT 25.805 198.815 25.975 198.985 ;
        RECT 57.335 199.325 57.505 199.495 ;
        RECT 56.665 197.615 56.835 197.785 ;
        RECT 45.635 191.825 45.805 191.995 ;
        RECT 46.095 191.825 46.265 191.995 ;
        RECT 46.555 191.825 46.725 191.995 ;
        RECT 47.015 191.825 47.185 191.995 ;
        RECT 47.475 191.825 47.645 191.995 ;
        RECT 48.865 191.845 49.035 192.015 ;
        RECT 44.665 190.465 44.835 190.635 ;
      LAYER met1 ;
        RECT 51.060 217.610 51.565 218.580 ;
        RECT 21.265 215.745 22.785 216.220 ;
        RECT 22.060 215.730 22.785 215.745 ;
        RECT 22.310 215.050 22.785 215.730 ;
        RECT 22.310 215.015 22.900 215.050 ;
        RECT 25.320 215.040 25.780 217.430 ;
        RECT 30.825 216.495 31.320 217.505 ;
        RECT 30.840 216.060 31.300 216.495 ;
        RECT 33.200 216.420 33.700 217.510 ;
        RECT 30.100 215.580 31.480 216.060 ;
        RECT 32.470 215.960 33.700 216.420 ;
        RECT 32.475 215.570 32.935 215.960 ;
        RECT 22.440 214.570 22.900 215.015 ;
        RECT 24.300 214.990 25.780 215.040 ;
        RECT 24.300 214.560 25.680 214.990 ;
        RECT 51.080 212.970 51.540 217.610 ;
        RECT 45.980 212.580 47.040 212.595 ;
        RECT 41.930 212.120 47.040 212.580 ;
        RECT 51.080 212.510 52.970 212.970 ;
        RECT 56.430 212.840 56.915 214.000 ;
        RECT 26.755 211.190 27.965 211.205 ;
        RECT 20.860 210.750 23.530 210.990 ;
        RECT 24.940 210.750 27.965 211.190 ;
        RECT 20.860 210.530 23.550 210.750 ;
        RECT 23.090 210.270 23.550 210.530 ;
        RECT 24.440 210.730 27.965 210.750 ;
        RECT 24.440 210.270 25.820 210.730 ;
        RECT 26.755 210.715 27.965 210.730 ;
        RECT 41.930 210.350 42.390 212.120 ;
        RECT 45.980 212.110 47.040 212.120 ;
        RECT 46.435 210.420 46.940 210.900 ;
        RECT 45.100 210.350 46.940 210.420 ;
        RECT 40.340 209.870 43.560 210.350 ;
        RECT 44.690 209.915 46.940 210.350 ;
        RECT 52.510 210.300 52.970 212.510 ;
        RECT 56.440 210.680 56.900 212.840 ;
        RECT 44.690 209.870 45.150 209.915 ;
        RECT 51.940 209.820 54.240 210.300 ;
        RECT 55.470 210.220 56.900 210.680 ;
        RECT 55.490 209.820 55.950 210.220 ;
        RECT 25.250 206.180 25.710 206.700 ;
        RECT 20.070 205.985 21.420 206.020 ;
        RECT 20.070 205.500 23.590 205.985 ;
        RECT 20.070 205.460 21.420 205.500 ;
        RECT 23.105 205.380 23.590 205.500 ;
        RECT 25.280 205.415 25.680 206.180 ;
        RECT 35.035 205.510 36.085 205.520 ;
        RECT 31.770 205.430 36.085 205.510 ;
        RECT 25.175 205.400 25.680 205.415 ;
        RECT 23.105 205.210 23.610 205.380 ;
        RECT 23.150 204.900 23.610 205.210 ;
        RECT 24.560 204.920 25.940 205.400 ;
        RECT 30.450 205.050 36.085 205.430 ;
        RECT 30.450 204.950 31.830 205.050 ;
        RECT 33.090 204.970 33.550 205.050 ;
        RECT 35.035 205.045 36.085 205.050 ;
        RECT 22.255 200.410 22.850 200.445 ;
        RECT 22.225 199.815 22.880 200.410 ;
        RECT 25.130 200.070 25.655 201.420 ;
        RECT 55.090 200.860 55.590 201.840 ;
        RECT 57.790 201.825 58.305 201.875 ;
        RECT 22.255 199.570 22.850 199.815 ;
        RECT 22.250 199.110 23.950 199.570 ;
        RECT 25.160 199.155 25.620 200.070 ;
        RECT 55.110 199.660 55.570 200.860 ;
        RECT 57.790 200.855 58.320 201.825 ;
        RECT 57.790 200.840 58.305 200.855 ;
        RECT 57.830 200.665 58.290 200.840 ;
        RECT 56.635 200.435 60.535 200.665 ;
        RECT 54.650 199.180 56.030 199.660 ;
        RECT 25.075 199.140 25.620 199.155 ;
        RECT 22.320 199.100 22.780 199.110 ;
        RECT 23.480 198.660 23.940 199.110 ;
        RECT 24.740 198.660 26.120 199.140 ;
        RECT 56.635 197.845 56.865 200.435 ;
        RECT 57.830 200.080 58.290 200.435 ;
        RECT 57.170 199.620 58.290 200.080 ;
        RECT 57.190 199.170 57.650 199.620 ;
        RECT 57.830 199.600 58.290 199.620 ;
        RECT 56.605 197.555 56.895 197.845 ;
        RECT 56.635 197.485 56.865 197.555 ;
        RECT 60.335 195.215 60.565 200.435 ;
        RECT 43.585 195.085 60.565 195.215 ;
        RECT 43.565 194.985 60.565 195.085 ;
        RECT 43.565 194.315 43.840 194.985 ;
        RECT 43.550 193.095 43.845 193.110 ;
        RECT 43.550 192.455 43.850 193.095 ;
        RECT 45.920 193.020 46.415 193.035 ;
        RECT 43.555 192.205 43.850 192.455 ;
        RECT 43.585 190.665 43.815 192.205 ;
        RECT 45.810 192.150 46.415 193.020 ;
        RECT 48.755 192.170 49.175 192.890 ;
        RECT 45.490 191.670 47.790 192.150 ;
        RECT 48.720 191.690 49.180 192.170 ;
        RECT 44.035 190.665 45.065 190.815 ;
        RECT 43.585 190.435 45.065 190.665 ;
        RECT 44.035 190.285 45.065 190.435 ;
      LAYER via ;
        RECT 51.170 218.190 51.430 218.450 ;
        RECT 25.420 217.000 25.680 217.260 ;
        RECT 21.520 215.850 21.780 216.110 ;
        RECT 30.940 217.070 31.200 217.330 ;
        RECT 33.320 217.020 33.580 217.280 ;
        RECT 56.540 213.460 56.800 213.720 ;
        RECT 46.550 212.220 46.810 212.480 ;
        RECT 21.000 210.630 21.260 210.890 ;
        RECT 27.330 210.830 27.590 211.090 ;
        RECT 46.550 210.490 46.810 210.750 ;
        RECT 25.350 206.310 25.610 206.570 ;
        RECT 20.490 205.560 20.750 205.820 ;
        RECT 35.600 205.150 35.860 205.410 ;
        RECT 55.210 201.440 55.470 201.700 ;
        RECT 25.260 200.880 25.520 201.140 ;
        RECT 22.260 199.820 22.840 200.400 ;
        RECT 57.930 201.440 58.190 201.700 ;
        RECT 43.570 194.370 43.830 194.630 ;
        RECT 43.570 192.570 43.830 192.830 ;
        RECT 46.020 192.610 46.280 192.870 ;
        RECT 48.840 192.580 49.100 192.840 ;
      LAYER met2 ;
        RECT 6.875 218.015 56.955 218.625 ;
        RECT 19.010 210.990 19.470 218.015 ;
        RECT 21.420 216.680 21.880 218.015 ;
        RECT 25.320 216.730 25.780 218.015 ;
        RECT 21.415 215.635 21.890 216.680 ;
        RECT 27.230 211.675 27.690 218.015 ;
        RECT 30.830 216.850 31.310 218.015 ;
        RECT 33.220 216.800 33.680 218.015 ;
        RECT 20.425 210.990 21.525 211.005 ;
        RECT 19.010 210.530 21.525 210.990 ;
        RECT 27.210 210.610 27.715 211.675 ;
        RECT 20.390 210.515 21.525 210.530 ;
        RECT 20.390 207.020 20.850 210.515 ;
        RECT 20.390 206.670 25.670 207.020 ;
        RECT 20.390 206.560 25.740 206.670 ;
        RECT 20.390 202.020 20.850 206.560 ;
        RECT 25.210 206.210 25.740 206.560 ;
        RECT 35.500 205.985 35.960 218.015 ;
        RECT 46.450 211.325 46.910 218.015 ;
        RECT 56.345 215.045 56.955 218.015 ;
        RECT 56.345 214.435 59.505 215.045 ;
        RECT 56.345 213.195 56.955 214.435 ;
        RECT 46.435 210.305 46.925 211.325 ;
        RECT 35.490 204.960 35.975 205.985 ;
        RECT 58.895 202.775 59.505 214.435 ;
        RECT 58.895 202.165 63.455 202.775 ;
        RECT 20.390 201.725 25.620 202.020 ;
        RECT 58.895 201.875 59.505 202.165 ;
        RECT 20.390 201.560 25.645 201.725 ;
        RECT 22.320 200.805 22.780 201.560 ;
        RECT 22.290 200.440 22.815 200.805 ;
        RECT 25.140 200.660 25.645 201.560 ;
        RECT 54.965 201.265 59.505 201.875 ;
        RECT 22.255 199.785 22.850 200.440 ;
        RECT 43.570 194.120 43.830 194.780 ;
        RECT 43.585 193.100 43.815 194.120 ;
        RECT 43.555 192.400 43.855 193.100 ;
        RECT 62.845 193.025 63.455 202.165 ;
        RECT 45.665 192.970 63.455 193.025 ;
        RECT 45.660 192.510 63.455 192.970 ;
        RECT 45.665 192.415 63.455 192.510 ;
      LAYER via2 ;
        RECT 7.110 218.180 7.390 218.460 ;
      LAYER met3 ;
        RECT 1.610 218.000 7.550 218.645 ;
      LAYER via3 ;
        RECT 1.705 218.160 2.025 218.480 ;
      LAYER met4 ;
        RECT 0.000 218.550 2.000 220.760 ;
        RECT 0.000 218.090 2.095 218.550 ;
        RECT 0.000 5.000 2.000 218.090 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 32.620 213.410 32.790 213.935 ;
        RECT 22.585 212.410 22.755 212.935 ;
        RECT 23.235 208.110 23.405 208.635 ;
        RECT 44.835 207.710 45.005 208.235 ;
        RECT 55.635 207.660 55.805 208.185 ;
        RECT 23.295 202.740 23.465 203.265 ;
        RECT 33.235 202.810 33.405 203.335 ;
        RECT 23.625 196.500 23.795 197.025 ;
        RECT 57.335 197.010 57.505 197.535 ;
        RECT 48.865 189.530 49.035 190.055 ;
      LAYER li1 ;
        RECT 30.205 213.185 30.445 213.995 ;
        RECT 31.115 213.185 31.385 213.995 ;
        RECT 30.100 213.015 31.480 213.185 ;
        RECT 32.560 213.175 32.850 213.900 ;
        RECT 32.475 213.005 32.935 213.175 ;
        RECT 22.525 212.175 22.815 212.900 ;
        RECT 22.440 212.005 22.900 212.175 ;
        RECT 24.620 212.165 24.850 212.985 ;
        RECT 24.300 211.995 25.680 212.165 ;
        RECT 23.775 209.105 24.025 209.110 ;
        RECT 23.775 208.865 25.090 209.105 ;
        RECT 53.915 208.870 54.155 209.295 ;
        RECT 23.775 208.860 24.025 208.865 ;
        RECT 23.175 207.875 23.465 208.600 ;
        RECT 24.760 207.875 24.990 208.695 ;
        RECT 41.180 208.465 41.730 208.665 ;
        RECT 53.915 208.630 54.920 208.870 ;
        RECT 53.915 208.315 54.155 208.630 ;
        RECT 23.090 207.705 23.550 207.875 ;
        RECT 24.440 207.705 25.820 207.875 ;
        RECT 40.475 207.475 40.805 207.865 ;
        RECT 41.315 207.475 41.645 207.865 ;
        RECT 43.185 207.475 43.475 208.310 ;
        RECT 44.775 207.475 45.065 208.200 ;
        RECT 40.340 207.305 43.560 207.475 ;
        RECT 44.690 207.305 45.150 207.475 ;
        RECT 52.455 207.425 53.390 207.825 ;
        RECT 55.575 207.425 55.865 208.150 ;
        RECT 51.940 207.255 54.240 207.425 ;
        RECT 55.490 207.255 55.950 207.425 ;
        RECT 30.545 204.725 30.875 204.920 ;
        RECT 29.625 204.555 30.875 204.725 ;
        RECT 30.545 204.135 30.875 204.555 ;
        RECT 30.545 203.965 31.225 204.135 ;
        RECT 23.895 203.795 24.225 203.800 ;
        RECT 23.820 203.755 24.540 203.795 ;
        RECT 23.820 203.515 25.210 203.755 ;
        RECT 23.820 203.475 24.540 203.515 ;
        RECT 23.895 203.470 24.225 203.475 ;
        RECT 31.055 203.365 31.225 203.965 ;
        RECT 23.235 202.505 23.525 203.230 ;
        RECT 24.880 202.525 25.110 203.345 ;
        RECT 30.555 202.555 30.795 203.365 ;
        RECT 30.965 202.725 31.295 203.365 ;
        RECT 31.465 202.555 31.735 203.365 ;
        RECT 33.175 202.575 33.465 203.300 ;
        RECT 23.150 202.335 23.610 202.505 ;
        RECT 24.560 202.355 25.940 202.525 ;
        RECT 30.450 202.385 31.830 202.555 ;
        RECT 33.090 202.405 33.550 202.575 ;
        RECT 23.565 196.265 23.855 196.990 ;
        RECT 25.060 196.265 25.290 197.085 ;
        RECT 54.970 196.785 55.200 197.605 ;
        RECT 54.650 196.615 56.030 196.785 ;
        RECT 57.275 196.775 57.565 197.500 ;
        RECT 57.190 196.605 57.650 196.775 ;
        RECT 23.480 196.095 23.940 196.265 ;
        RECT 24.740 196.095 26.120 196.265 ;
        RECT 47.110 191.315 47.705 191.655 ;
        RECT 47.110 189.995 47.285 191.315 ;
        RECT 47.465 190.720 47.705 191.145 ;
        RECT 47.465 190.480 48.350 190.720 ;
        RECT 47.465 190.165 47.705 190.480 ;
        RECT 47.110 189.825 47.705 189.995 ;
        RECT 46.005 189.275 46.940 189.675 ;
        RECT 47.110 189.655 48.485 189.825 ;
        RECT 47.110 189.445 47.705 189.655 ;
        RECT 48.805 189.295 49.095 190.020 ;
        RECT 45.490 189.105 47.790 189.275 ;
        RECT 48.720 189.125 49.180 189.295 ;
      LAYER mcon ;
        RECT 30.245 213.015 30.415 213.185 ;
        RECT 30.705 213.015 30.875 213.185 ;
        RECT 31.165 213.015 31.335 213.185 ;
        RECT 32.620 213.005 32.790 213.175 ;
        RECT 22.585 212.005 22.755 212.175 ;
        RECT 24.445 211.995 24.615 212.165 ;
        RECT 24.905 211.995 25.075 212.165 ;
        RECT 25.365 211.995 25.535 212.165 ;
        RECT 23.815 208.900 23.985 209.070 ;
        RECT 41.365 208.465 41.535 208.635 ;
        RECT 54.715 208.660 54.885 208.830 ;
        RECT 23.235 207.705 23.405 207.875 ;
        RECT 24.585 207.705 24.755 207.875 ;
        RECT 25.045 207.705 25.215 207.875 ;
        RECT 25.505 207.705 25.675 207.875 ;
        RECT 40.485 207.305 40.655 207.475 ;
        RECT 40.945 207.305 41.115 207.475 ;
        RECT 41.405 207.305 41.575 207.475 ;
        RECT 41.865 207.305 42.035 207.475 ;
        RECT 42.325 207.305 42.495 207.475 ;
        RECT 42.785 207.305 42.955 207.475 ;
        RECT 43.245 207.305 43.415 207.475 ;
        RECT 44.835 207.305 45.005 207.475 ;
        RECT 52.085 207.255 52.255 207.425 ;
        RECT 52.545 207.255 52.715 207.425 ;
        RECT 53.005 207.255 53.175 207.425 ;
        RECT 53.465 207.255 53.635 207.425 ;
        RECT 53.925 207.255 54.095 207.425 ;
        RECT 55.635 207.255 55.805 207.425 ;
        RECT 23.975 203.550 24.145 203.720 ;
        RECT 23.295 202.335 23.465 202.505 ;
        RECT 24.705 202.355 24.875 202.525 ;
        RECT 25.165 202.355 25.335 202.525 ;
        RECT 25.625 202.355 25.795 202.525 ;
        RECT 30.595 202.385 30.765 202.555 ;
        RECT 31.055 202.385 31.225 202.555 ;
        RECT 31.515 202.385 31.685 202.555 ;
        RECT 33.235 202.405 33.405 202.575 ;
        RECT 54.795 196.615 54.965 196.785 ;
        RECT 55.255 196.615 55.425 196.785 ;
        RECT 55.715 196.615 55.885 196.785 ;
        RECT 57.335 196.605 57.505 196.775 ;
        RECT 23.625 196.095 23.795 196.265 ;
        RECT 24.885 196.095 25.055 196.265 ;
        RECT 25.345 196.095 25.515 196.265 ;
        RECT 25.805 196.095 25.975 196.265 ;
        RECT 48.095 190.515 48.265 190.685 ;
        RECT 48.315 189.655 48.485 189.825 ;
        RECT 45.635 189.105 45.805 189.275 ;
        RECT 46.095 189.105 46.265 189.275 ;
        RECT 46.555 189.105 46.725 189.275 ;
        RECT 47.015 189.105 47.185 189.275 ;
        RECT 47.475 189.105 47.645 189.275 ;
        RECT 48.865 189.125 49.035 189.295 ;
      LAYER met1 ;
        RECT 30.100 212.955 31.480 213.340 ;
        RECT 32.475 212.955 32.935 213.330 ;
        RECT 30.100 212.910 32.935 212.955 ;
        RECT 30.050 212.850 32.935 212.910 ;
        RECT 30.050 212.800 32.925 212.850 ;
        RECT 7.145 211.995 7.465 212.050 ;
        RECT 22.440 211.995 22.900 212.330 ;
        RECT 24.300 211.995 25.680 212.320 ;
        RECT 7.145 211.840 25.680 211.995 ;
        RECT 7.145 211.790 7.465 211.840 ;
        RECT 19.815 211.255 24.025 211.505 ;
        RECT 12.040 210.425 12.910 210.460 ;
        RECT 19.815 210.425 20.065 211.255 ;
        RECT 23.775 210.970 24.025 211.255 ;
        RECT 12.040 210.175 20.075 210.425 ;
        RECT 12.040 210.140 12.910 210.175 ;
        RECT 23.775 209.170 24.285 210.970 ;
        RECT 23.745 208.800 24.285 209.170 ;
        RECT 23.090 207.625 23.550 208.030 ;
        RECT 23.075 207.550 23.550 207.625 ;
        RECT 23.075 207.465 23.325 207.550 ;
        RECT 8.460 207.345 23.325 207.465 ;
        RECT 23.880 207.345 24.285 208.800 ;
        RECT 24.440 207.550 25.820 208.030 ;
        RECT 24.615 207.345 24.770 207.550 ;
        RECT 30.050 207.345 30.425 212.800 ;
        RECT 41.315 208.365 41.635 208.735 ;
        RECT 54.630 208.625 55.225 208.870 ;
        RECT 8.460 207.140 30.425 207.345 ;
        RECT 8.475 206.985 30.425 207.140 ;
        RECT 38.665 207.985 38.835 208.000 ;
        RECT 41.365 207.985 41.535 208.365 ;
        RECT 38.665 207.815 41.535 207.985 ;
        RECT 9.450 206.965 23.320 206.985 ;
        RECT 12.110 203.660 12.495 204.345 ;
        RECT 12.165 203.565 12.435 203.660 ;
        RECT 12.215 187.435 12.385 203.565 ;
        RECT 15.900 202.355 16.400 206.965 ;
        RECT 23.880 206.615 24.285 206.985 ;
        RECT 19.430 206.285 24.285 206.615 ;
        RECT 19.430 205.285 19.760 206.285 ;
        RECT 19.430 204.930 19.765 205.285 ;
        RECT 19.425 204.530 19.765 204.930 ;
        RECT 23.880 203.830 24.285 206.285 ;
        RECT 38.665 206.185 38.835 207.815 ;
        RECT 40.340 207.150 43.560 207.630 ;
        RECT 44.690 207.150 45.150 207.630 ;
        RECT 28.985 206.015 38.835 206.185 ;
        RECT 28.985 204.725 29.155 206.015 ;
        RECT 38.665 205.250 38.835 206.015 ;
        RECT 41.985 206.575 42.275 207.150 ;
        RECT 44.825 206.575 44.980 207.150 ;
        RECT 51.940 207.100 54.240 207.580 ;
        RECT 53.635 206.575 53.920 207.100 ;
        RECT 41.985 206.275 53.920 206.575 ;
        RECT 40.950 205.250 41.600 205.400 ;
        RECT 38.650 205.050 41.700 205.250 ;
        RECT 29.595 204.725 29.825 204.785 ;
        RECT 28.985 204.555 29.975 204.725 ;
        RECT 29.595 204.495 29.825 204.555 ;
        RECT 23.865 203.440 24.285 203.830 ;
        RECT 23.880 203.390 24.285 203.440 ;
        RECT 23.150 202.355 23.610 202.660 ;
        RECT 24.560 202.385 25.940 202.680 ;
        RECT 30.450 202.385 31.830 202.710 ;
        RECT 24.560 202.355 31.830 202.385 ;
        RECT 15.900 202.230 31.830 202.355 ;
        RECT 33.090 202.250 33.550 202.730 ;
        RECT 15.900 202.200 25.940 202.230 ;
        RECT 15.900 196.100 16.400 202.200 ;
        RECT 23.150 202.180 23.610 202.200 ;
        RECT 23.480 196.100 23.940 196.420 ;
        RECT 24.740 196.100 26.120 196.420 ;
        RECT 33.240 196.100 33.395 202.250 ;
        RECT 38.650 197.655 38.850 205.050 ;
        RECT 40.950 204.900 41.600 205.050 ;
        RECT 41.985 204.480 42.275 206.275 ;
        RECT 42.590 205.250 42.910 205.280 ;
        RECT 54.980 205.250 55.225 208.625 ;
        RECT 55.490 207.100 55.950 207.580 ;
        RECT 42.590 205.080 55.225 205.250 ;
        RECT 42.590 205.050 55.200 205.080 ;
        RECT 42.590 205.020 42.910 205.050 ;
        RECT 55.625 204.480 55.780 207.100 ;
        RECT 41.985 204.325 55.775 204.480 ;
        RECT 38.600 196.850 38.905 197.655 ;
        RECT 38.650 196.100 38.850 196.850 ;
        RECT 41.985 196.615 42.275 204.325 ;
        RECT 54.650 196.655 56.030 196.940 ;
        RECT 57.190 196.655 57.650 196.930 ;
        RECT 54.650 196.615 57.655 196.655 ;
        RECT 41.985 196.460 57.655 196.615 ;
        RECT 41.985 196.100 42.275 196.460 ;
        RECT 57.190 196.450 57.650 196.460 ;
        RECT 15.900 195.605 42.275 196.100 ;
        RECT 15.900 195.600 42.250 195.605 ;
        RECT 36.575 189.105 36.730 195.600 ;
        RECT 38.650 195.370 38.850 195.600 ;
        RECT 38.630 195.240 38.870 195.370 ;
        RECT 38.610 194.460 38.895 195.240 ;
        RECT 38.650 193.550 38.850 194.460 ;
        RECT 38.650 193.350 48.320 193.550 ;
        RECT 38.650 189.105 38.850 193.350 ;
        RECT 48.110 190.720 48.310 193.350 ;
        RECT 48.030 190.700 48.330 190.720 ;
        RECT 48.030 190.500 48.390 190.700 ;
        RECT 48.030 190.480 48.330 190.500 ;
        RECT 48.280 189.460 48.520 189.890 ;
        RECT 45.490 189.105 47.790 189.430 ;
        RECT 36.575 188.950 47.825 189.105 ;
        RECT 47.275 188.330 47.430 188.950 ;
        RECT 47.570 188.330 47.830 188.410 ;
        RECT 47.275 188.175 47.830 188.330 ;
        RECT 47.570 188.090 47.830 188.175 ;
        RECT 48.315 187.435 48.485 189.460 ;
        RECT 48.720 189.130 49.180 189.450 ;
        RECT 48.720 188.970 49.890 189.130 ;
        RECT 48.945 188.950 49.890 188.970 ;
        RECT 48.950 188.830 49.890 188.950 ;
        RECT 49.590 188.400 49.890 188.830 ;
        RECT 48.800 188.100 49.890 188.400 ;
        RECT 12.215 187.265 48.485 187.435 ;
      LAYER via ;
        RECT 7.175 211.790 7.435 212.050 ;
        RECT 12.170 210.170 12.430 210.430 ;
        RECT 8.670 207.095 8.930 207.355 ;
        RECT 12.170 203.920 12.430 204.180 ;
        RECT 19.470 204.670 19.730 204.930 ;
        RECT 41.170 205.020 41.430 205.280 ;
        RECT 42.620 205.020 42.880 205.280 ;
        RECT 38.620 197.020 38.880 197.280 ;
        RECT 38.625 194.920 38.885 195.180 ;
        RECT 47.570 188.120 47.830 188.380 ;
        RECT 48.975 188.125 49.235 188.385 ;
      LAYER met2 ;
        RECT 6.030 212.050 6.470 212.100 ;
        RECT 7.175 212.050 7.435 212.080 ;
        RECT 6.030 211.800 7.435 212.050 ;
        RECT 6.030 211.750 6.470 211.800 ;
        RECT 7.175 211.760 7.435 211.800 ;
        RECT 12.175 210.515 12.425 210.575 ;
        RECT 12.135 210.170 12.470 210.515 ;
        RECT 7.460 206.985 9.140 207.465 ;
        RECT 12.175 204.925 12.425 210.170 ;
        RECT 41.100 205.250 41.650 205.400 ;
        RECT 42.620 205.250 42.880 205.310 ;
        RECT 41.100 205.050 43.150 205.250 ;
        RECT 19.135 204.940 19.795 204.995 ;
        RECT 19.135 204.925 19.815 204.940 ;
        RECT 12.175 204.920 19.815 204.925 ;
        RECT 12.080 204.675 19.815 204.920 ;
        RECT 41.100 204.900 41.650 205.050 ;
        RECT 42.620 204.990 42.880 205.050 ;
        RECT 12.080 203.780 12.525 204.675 ;
        RECT 19.135 204.605 19.815 204.675 ;
        RECT 12.120 203.770 12.485 203.780 ;
        RECT 38.595 196.895 38.905 197.405 ;
        RECT 38.650 195.475 38.850 196.895 ;
        RECT 38.630 195.445 38.875 195.475 ;
        RECT 38.610 194.710 38.895 195.445 ;
        RECT 47.540 188.365 49.460 188.410 ;
        RECT 47.540 188.120 49.475 188.365 ;
        RECT 47.615 188.110 49.475 188.120 ;
      LAYER via2 ;
        RECT 6.110 211.785 6.390 212.065 ;
        RECT 7.610 207.085 7.890 207.365 ;
      LAYER met3 ;
        RECT 4.945 212.100 5.455 212.150 ;
        RECT 6.050 212.100 6.450 212.125 ;
        RECT 4.945 211.750 6.450 212.100 ;
        RECT 4.945 211.700 5.455 211.750 ;
        RECT 6.050 211.725 6.450 211.750 ;
        RECT 7.485 207.465 8.015 207.490 ;
        RECT 6.210 206.985 8.015 207.465 ;
        RECT 7.485 206.960 8.015 206.985 ;
      LAYER via3 ;
        RECT 5.040 211.765 5.360 212.085 ;
        RECT 6.490 207.065 6.810 207.385 ;
      LAYER met4 ;
        RECT 3.000 212.155 5.000 220.760 ;
        RECT 3.000 211.695 5.430 212.155 ;
        RECT 3.000 207.465 5.000 211.695 ;
        RECT 6.405 207.465 6.895 207.470 ;
        RECT 3.000 206.985 6.895 207.465 ;
        RECT 3.000 5.000 5.000 206.985 ;
        RECT 6.405 206.980 6.895 206.985 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 30.250 213.015 30.420 213.185 ;
        RECT 24.445 211.995 24.615 212.165 ;
        RECT 24.585 207.705 24.755 207.875 ;
        RECT 40.485 207.305 40.655 207.475 ;
        RECT 52.090 207.255 52.260 207.425 ;
        RECT 24.705 202.355 24.875 202.525 ;
        RECT 30.600 202.385 30.770 202.555 ;
        RECT 54.795 196.615 54.965 196.785 ;
        RECT 24.885 196.095 25.055 196.265 ;
        RECT 45.640 189.105 45.810 189.275 ;
      LAYER li1 ;
        RECT 30.195 215.355 30.525 215.550 ;
        RECT 29.465 215.185 30.525 215.355 ;
        RECT 30.195 214.765 30.525 215.185 ;
        RECT 30.195 214.595 30.875 214.765 ;
        RECT 25.020 213.565 25.350 214.545 ;
        RECT 29.075 214.175 30.535 214.425 ;
        RECT 30.705 213.995 30.875 214.595 ;
        RECT 31.045 214.175 32.245 214.425 ;
        RECT 25.120 213.215 25.350 213.565 ;
        RECT 30.615 213.355 30.945 213.995 ;
        RECT 25.120 212.985 26.515 213.215 ;
        RECT 25.120 212.965 25.350 212.985 ;
        RECT 25.020 212.335 25.350 212.965 ;
        RECT 25.160 209.275 25.490 210.255 ;
        RECT 25.260 208.915 25.490 209.275 ;
        RECT 40.425 209.175 40.805 209.855 ;
        RECT 41.735 209.345 42.065 209.855 ;
        RECT 42.575 209.345 42.975 209.855 ;
        RECT 41.735 209.175 42.975 209.345 ;
        RECT 43.155 209.265 43.475 209.855 ;
        RECT 52.025 209.405 52.285 209.805 ;
        RECT 25.260 208.685 26.615 208.915 ;
        RECT 25.260 208.675 25.490 208.685 ;
        RECT 25.160 208.045 25.490 208.675 ;
        RECT 40.425 208.215 40.595 209.175 ;
        RECT 43.155 209.095 44.385 209.265 ;
        RECT 52.025 209.235 53.390 209.405 ;
        RECT 40.765 208.835 42.070 209.005 ;
        RECT 43.155 208.925 43.475 209.095 ;
        RECT 52.025 209.045 52.485 209.065 ;
        RECT 50.520 209.015 52.485 209.045 ;
        RECT 40.765 208.385 41.010 208.835 ;
        RECT 41.900 208.635 42.070 208.835 ;
        RECT 42.845 208.755 43.475 208.925 ;
        RECT 41.900 208.465 42.275 208.635 ;
        RECT 42.445 208.215 42.675 208.715 ;
        RECT 40.425 208.045 42.675 208.215 ;
        RECT 40.975 207.725 41.145 208.045 ;
        RECT 42.845 207.875 43.015 208.755 ;
        RECT 50.500 208.615 52.485 209.015 ;
        RECT 50.520 208.585 52.485 208.615 ;
        RECT 52.025 208.335 52.485 208.585 ;
        RECT 52.655 208.165 53.390 209.235 ;
        RECT 42.060 207.705 43.015 207.875 ;
        RECT 52.025 207.995 53.390 208.165 ;
        RECT 52.025 207.595 52.285 207.995 ;
        RECT 25.280 203.925 25.610 204.905 ;
        RECT 25.380 203.615 25.610 203.925 ;
        RECT 30.535 203.790 30.885 203.795 ;
        RECT 25.380 203.385 27.085 203.615 ;
        RECT 29.600 203.545 30.885 203.790 ;
        RECT 31.395 203.545 32.645 203.795 ;
        RECT 25.380 203.325 25.610 203.385 ;
        RECT 25.280 202.695 25.610 203.325 ;
        RECT 25.460 197.665 25.790 198.645 ;
        RECT 54.180 197.775 55.300 198.015 ;
        RECT 25.560 197.315 25.790 197.665 ;
        RECT 25.560 197.085 27.015 197.315 ;
        RECT 25.560 197.065 25.790 197.085 ;
        RECT 25.460 196.435 25.790 197.065 ;
        RECT 45.575 191.255 45.835 191.655 ;
        RECT 45.575 191.085 46.940 191.255 ;
        RECT 46.205 190.015 46.940 191.085 ;
        RECT 45.575 189.845 46.940 190.015 ;
        RECT 45.575 189.445 45.835 189.845 ;
      LAYER mcon ;
        RECT 29.115 214.215 29.285 214.385 ;
        RECT 31.995 214.215 32.165 214.385 ;
        RECT 26.265 213.015 26.435 213.185 ;
        RECT 26.415 208.715 26.585 208.885 ;
        RECT 44.215 209.095 44.385 209.265 ;
        RECT 40.765 208.815 40.935 208.985 ;
        RECT 50.615 208.730 50.785 208.900 ;
        RECT 26.885 203.415 27.055 203.585 ;
        RECT 29.675 203.580 29.845 203.750 ;
        RECT 32.445 203.585 32.615 203.755 ;
        RECT 54.265 197.810 54.435 197.980 ;
        RECT 26.805 197.115 26.975 197.285 ;
      LAYER met1 ;
        RECT 159.180 218.620 161.000 219.060 ;
        RECT 26.675 217.890 32.205 217.895 ;
        RECT 26.675 217.645 32.240 217.890 ;
        RECT 26.685 213.215 26.915 217.645 ;
        RECT 29.405 215.355 29.695 215.385 ;
        RECT 28.765 215.185 29.695 215.355 ;
        RECT 28.765 215.030 28.935 215.185 ;
        RECT 29.405 215.155 29.695 215.185 ;
        RECT 28.690 214.770 29.010 215.030 ;
        RECT 31.960 214.425 32.240 217.645 ;
        RECT 26.185 212.985 26.915 213.215 ;
        RECT 28.525 214.175 29.355 214.425 ;
        RECT 31.915 214.175 32.275 214.425 ;
        RECT 28.525 208.915 28.775 214.175 ;
        RECT 31.960 214.160 32.240 214.175 ;
        RECT 30.940 212.385 31.260 212.430 ;
        RECT 30.940 212.215 38.935 212.385 ;
        RECT 30.940 212.170 31.260 212.215 ;
        RECT 26.355 208.685 28.775 208.915 ;
        RECT 38.765 208.985 38.935 212.215 ;
        RECT 44.215 211.215 50.035 211.235 ;
        RECT 44.185 211.065 50.035 211.215 ;
        RECT 44.185 209.265 44.420 211.065 ;
        RECT 44.115 209.095 44.420 209.265 ;
        RECT 40.665 208.985 41.035 209.085 ;
        RECT 44.185 209.035 44.420 209.095 ;
        RECT 49.570 209.045 50.035 211.065 ;
        RECT 38.765 208.815 41.035 208.985 ;
        RECT 40.665 208.715 41.035 208.815 ;
        RECT 49.570 208.585 50.980 209.045 ;
        RECT 49.580 207.060 49.820 208.585 ;
        RECT 49.570 206.740 49.830 207.060 ;
        RECT 29.640 203.790 29.885 203.820 ;
        RECT 26.825 203.615 27.115 203.645 ;
        RECT 27.410 203.615 30.020 203.790 ;
        RECT 26.765 203.545 30.020 203.615 ;
        RECT 26.765 203.385 27.645 203.545 ;
        RECT 29.640 203.515 29.885 203.545 ;
        RECT 26.825 203.355 27.115 203.385 ;
        RECT 32.330 203.180 32.670 203.820 ;
        RECT 49.570 203.270 49.830 203.730 ;
        RECT 26.745 197.315 27.035 197.345 ;
        RECT 32.360 197.315 32.640 203.180 ;
        RECT 49.430 202.780 49.920 203.270 ;
        RECT 49.580 198.015 49.820 202.780 ;
        RECT 49.580 197.775 54.520 198.015 ;
        RECT 26.705 197.085 32.635 197.315 ;
        RECT 26.745 197.055 27.035 197.085 ;
      LAYER via ;
        RECT 28.720 214.770 28.980 215.030 ;
        RECT 30.970 212.170 31.230 212.430 ;
        RECT 49.570 206.770 49.830 207.030 ;
        RECT 49.570 203.020 49.830 203.280 ;
      LAYER met2 ;
        RECT 28.720 214.740 28.980 215.060 ;
        RECT 28.765 212.385 28.935 214.740 ;
        RECT 30.970 212.385 31.230 212.460 ;
        RECT 28.765 212.215 31.230 212.385 ;
        RECT 30.970 212.140 31.230 212.215 ;
        RECT 49.540 207.025 49.860 207.030 ;
        RECT 49.455 206.770 49.860 207.025 ;
        RECT 49.455 203.520 49.845 206.770 ;
        RECT 49.430 202.880 49.920 203.520 ;
  END
END tt_um_template
END LIBRARY

