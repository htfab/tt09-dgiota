VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_17
  CLASS BLOCK ;
  FOREIGN tt_um_test_17 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 142.860 224.760 143.160 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 145.620 224.760 145.920 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 140.100 224.760 140.400 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 150.840 0.000 151.740 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 131.520 0.000 132.420 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 112.200 0.000 113.100 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 92.880 0.000 93.780 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 73.560 0.000 74.460 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 54.240 0.000 55.140 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 34.920 0.000 35.820 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 15.600 0.000 16.500 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 137.340 224.760 137.640 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 134.580 224.760 134.880 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 131.820 224.760 132.120 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 129.060 224.760 129.360 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 126.300 224.760 126.600 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 123.540 224.760 123.840 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 120.780 224.760 121.080 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 118.020 224.760 118.320 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 115.260 224.760 115.560 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 112.500 224.760 112.800 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 109.740 224.760 110.040 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 106.980 224.760 107.280 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 104.220 224.760 104.520 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 101.460 224.760 101.760 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 98.700 224.760 99.000 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 95.940 224.760 96.240 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 49.020 224.760 49.320 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 46.260 224.760 46.560 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 43.500 224.760 43.800 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 40.740 224.760 41.040 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 37.980 224.760 38.280 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 35.220 224.760 35.520 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 32.460 224.760 32.760 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 29.700 224.760 30.000 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 71.100 224.760 71.400 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 68.340 224.760 68.640 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 65.580 224.760 65.880 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 62.820 224.760 63.120 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 60.060 224.760 60.360 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 57.300 224.760 57.600 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 54.540 224.760 54.840 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 51.780 224.760 52.080 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 93.180 224.760 93.480 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 90.420 224.760 90.720 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 87.660 224.760 87.960 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 84.900 224.760 85.200 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 82.140 224.760 82.440 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 79.380 224.760 79.680 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 76.620 224.760 76.920 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 73.860 224.760 74.160 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.030 5.000 2.030 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.030 5.000 5.030 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 22.190 140.315 56.570 175.460 ;
      LAYER li1 ;
        RECT 21.630 140.305 56.380 175.355 ;
      LAYER met1 ;
        RECT 13.780 131.250 161.000 225.750 ;
      LAYER met2 ;
        RECT 17.980 73.565 118.730 176.885 ;
      LAYER met3 ;
        RECT 0.000 0.020 151.730 179.400 ;
      LAYER met4 ;
        RECT 2.430 4.600 2.630 171.055 ;
        RECT 5.430 4.600 150.840 171.055 ;
        RECT 0.025 1.400 150.840 4.600 ;
        RECT 0.025 0.045 15.200 1.400 ;
        RECT 16.900 0.045 34.520 1.400 ;
        RECT 36.220 0.045 53.840 1.400 ;
        RECT 55.540 0.045 73.160 1.400 ;
        RECT 74.860 0.045 92.480 1.400 ;
        RECT 94.180 0.045 111.800 1.400 ;
        RECT 113.500 0.045 131.120 1.400 ;
        RECT 132.820 0.045 150.440 1.400 ;
  END
END tt_um_test_17
END LIBRARY

