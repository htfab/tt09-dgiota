magic
tech sky130A
magscale 1 2
timestamp 1731205162
<< nwell >>
rect 6139 35090 6716 35092
rect 6139 34771 7064 35090
rect 6712 34769 7064 34771
rect 7659 34432 8236 34492
rect 7659 34171 8586 34432
rect 8232 34111 8586 34171
rect 6049 34030 6536 34032
rect 6049 33711 6844 34030
rect 6532 33709 6844 33711
rect 10305 32760 10886 32770
rect 10305 32449 11244 32760
rect 10872 32439 11244 32449
rect 6332 32262 6674 32270
rect 5839 31949 6674 32262
rect 5839 31941 6356 31949
rect 7809 31760 8386 31762
rect 7809 31441 8724 31760
rect 8382 31439 8724 31441
rect 5847 30969 6644 31290
rect 7327 29070 7816 29080
rect 5312 29032 5644 29040
rect 4653 28719 5644 29032
rect 7327 28759 8114 29070
rect 7782 28749 8114 28759
rect 4653 28711 5316 28719
rect 10363 28660 10966 28662
rect 10363 28341 11314 28660
rect 10962 28339 11314 28341
<< locali >>
rect 6006 34767 6238 34770
rect 6006 34733 6009 34767
rect 6043 34733 6238 34767
rect 6006 34730 6238 34733
rect 6310 34737 6629 34743
rect 6310 34703 6589 34737
rect 6623 34703 6629 34737
rect 6310 34697 6629 34703
rect 7536 34617 7666 34620
rect 7536 34583 7619 34617
rect 7653 34583 7666 34617
rect 7536 34580 7666 34583
rect 7536 34350 7576 34580
rect 7536 34310 7746 34350
rect 7896 34167 8165 34169
rect 7896 34133 8129 34167
rect 8163 34133 8165 34167
rect 7896 34131 8165 34133
rect 5896 33707 6148 33710
rect 5896 33673 5899 33707
rect 5933 33673 6148 33707
rect 5896 33670 6148 33673
rect 6220 33677 6519 33683
rect 6220 33643 6479 33677
rect 6513 33643 6519 33677
rect 6220 33637 6519 33643
rect 10537 32550 10571 32563
rect 10537 32540 10586 32550
rect 10574 32500 10586 32540
rect 10566 32490 10586 32500
rect 10029 32449 10078 32486
rect 10063 32415 10078 32449
rect 10029 32406 10078 32415
rect 10146 32409 10213 32443
rect 5676 31937 5938 31940
rect 5676 31903 5679 31937
rect 5713 31903 5938 31937
rect 5676 31900 5938 31903
rect 6010 31877 6319 31903
rect 6010 31857 6279 31877
rect 6273 31843 6279 31857
rect 6313 31843 6319 31877
rect 6273 31827 6319 31843
rect 7806 31610 7836 31620
rect 7806 31570 7823 31610
rect 7806 31560 7836 31570
rect 7621 31439 7853 31445
rect 7621 31401 7657 31439
rect 7695 31401 7853 31439
rect 7946 31412 7962 31460
rect 8032 31440 8048 31445
rect 8032 31437 8266 31440
rect 8032 31403 8219 31437
rect 8253 31403 8266 31437
rect 8032 31402 8266 31403
rect 7621 31395 7853 31401
rect 8045 31400 8266 31402
rect 5686 30967 5946 30970
rect 5686 30933 5689 30967
rect 5723 30933 5946 30967
rect 6273 30958 6319 30983
rect 6273 30933 6278 30958
rect 5686 30930 5946 30933
rect 6018 30922 6278 30933
rect 6314 30922 6319 30958
rect 6018 30887 6319 30922
rect 7216 28720 7406 28760
rect 4326 28697 4523 28700
rect 4326 28663 4329 28697
rect 4363 28663 4523 28697
rect 4326 28660 4523 28663
rect 4892 28687 5106 28690
rect 4892 28653 5069 28687
rect 5103 28653 5106 28687
rect 4892 28650 5106 28653
rect 10026 28329 10206 28330
rect 10026 28327 10233 28329
rect 10026 28293 10029 28327
rect 10063 28293 10233 28327
rect 10026 28290 10233 28293
rect 10602 28327 10846 28330
rect 10602 28293 10809 28327
rect 10843 28293 10846 28327
rect 10602 28290 10846 28293
rect 10582 28214 10786 28220
rect 10582 28166 10732 28214
rect 10780 28166 10786 28214
rect 10582 28160 10786 28166
<< viali >>
rect 6009 34733 6043 34767
rect 6589 34703 6623 34737
rect 7619 34583 7653 34617
rect 7709 34133 7743 34167
rect 8129 34133 8163 34167
rect 5899 33673 5933 33707
rect 6479 33643 6513 33677
rect 10534 32500 10574 32540
rect 10029 32415 10063 32449
rect 10112 32409 10146 32443
rect 5679 31903 5713 31937
rect 6279 31843 6313 31877
rect 7823 31570 7863 31610
rect 7657 31401 7695 31439
rect 8219 31403 8253 31437
rect 5689 30933 5723 30967
rect 6278 30922 6314 30958
rect 7176 28720 7216 28760
rect 7499 28703 7533 28737
rect 4329 28663 4363 28697
rect 5069 28653 5103 28687
rect 4879 28543 4913 28577
rect 10029 28293 10063 28327
rect 10809 28293 10843 28327
rect 10732 28166 10780 28214
<< metal1 >>
rect 29820 45090 32200 45150
rect 29820 45080 29880 45090
rect 6583 35657 7479 35703
rect 6298 35280 6356 35286
rect 6356 35220 6359 35279
rect 6298 35214 6359 35220
rect 6301 35044 6359 35214
rect 5997 34770 6055 34773
rect 2756 34767 6055 34770
rect 2756 34733 6009 34767
rect 6043 34733 6055 34767
rect 2756 34730 6055 34733
rect 2756 26310 2816 34730
rect 5997 34727 6055 34730
rect 6583 34737 6629 35657
rect 6946 35370 7006 35376
rect 6946 35054 7006 35310
rect 6583 34703 6589 34737
rect 6623 34703 6629 34737
rect 6583 34691 6629 34703
rect 4778 34410 4836 34416
rect 4777 34351 4778 34409
rect 6209 34409 6267 34520
rect 4836 34351 6267 34409
rect 6956 34420 7016 34505
rect 6956 34354 7016 34360
rect 4778 34344 4836 34350
rect 6473 34237 7279 34283
rect 5647 34131 6177 34189
rect 4788 34040 4846 34046
rect 4787 33981 4788 34039
rect 5647 34039 5705 34131
rect 4846 33981 5705 34039
rect 6119 33984 6177 34131
rect 4788 33974 4846 33980
rect 5887 33710 5945 33713
rect 4896 33707 5945 33710
rect 4896 33673 5899 33707
rect 5933 33673 5945 33707
rect 4896 33670 5945 33673
rect 4700 31946 4752 31952
rect 3396 31900 4700 31940
rect 3396 27100 3456 31900
rect 4700 31888 4752 31894
rect 4896 30970 4936 33670
rect 5887 33667 5945 33670
rect 6473 33677 6519 34237
rect 6726 34170 6785 34176
rect 6726 33995 6785 34110
rect 7233 33733 7279 34237
rect 7433 34173 7479 35657
rect 8016 34780 8926 34820
rect 7607 34620 7665 34623
rect 8016 34620 8056 34780
rect 8476 34660 8536 34666
rect 7606 34617 8056 34620
rect 7606 34583 7619 34617
rect 7653 34583 8056 34617
rect 7606 34580 8056 34583
rect 8475 34600 8476 34660
rect 8475 34594 8536 34600
rect 7607 34577 7665 34580
rect 8026 34480 8086 34486
rect 7936 34420 8026 34480
rect 8026 34414 8086 34420
rect 8475 34396 8535 34594
rect 7433 34167 7755 34173
rect 7433 34133 7709 34167
rect 7743 34133 7755 34167
rect 7433 34127 7755 34133
rect 8123 34167 8169 34179
rect 8123 34133 8129 34167
rect 8163 34133 8169 34167
rect 7538 33920 7596 33926
rect 7537 33862 7538 33920
rect 7596 33862 7787 33920
rect 7538 33854 7596 33860
rect 8123 33733 8169 34133
rect 7233 33687 8169 33733
rect 8466 33720 8526 33847
rect 6473 33643 6479 33677
rect 6513 33643 6519 33677
rect 8466 33654 8526 33660
rect 6473 33631 6519 33643
rect 5138 33300 5196 33306
rect 5137 33241 5138 33299
rect 6119 33299 6177 33460
rect 5196 33241 6177 33299
rect 6725 33336 6785 33445
rect 6725 33330 6786 33336
rect 6725 33270 6726 33330
rect 6726 33264 6786 33270
rect 5138 33234 5196 33240
rect 6273 32507 7539 32553
rect 5908 32470 5966 32476
rect 5966 32410 5967 32469
rect 5908 32404 5967 32410
rect 5909 32214 5967 32404
rect 5120 31946 5172 31952
rect 5667 31940 5725 31943
rect 5172 31937 5725 31940
rect 5172 31903 5679 31937
rect 5713 31903 5725 31937
rect 5172 31900 5725 31903
rect 5667 31897 5725 31900
rect 5120 31888 5172 31894
rect 6273 31877 6319 32507
rect 6726 32430 6785 32436
rect 6556 32370 6726 32429
rect 6556 32235 6615 32370
rect 6726 32364 6785 32370
rect 6273 31843 6279 31877
rect 6313 31843 6319 31877
rect 6273 31831 6319 31843
rect 5118 31570 5176 31576
rect 5117 31511 5118 31569
rect 5909 31569 5967 31690
rect 6555 31650 6615 31685
rect 6726 31650 6786 31656
rect 6555 31590 6726 31650
rect 6726 31584 6786 31590
rect 5176 31511 5967 31569
rect 5118 31504 5176 31510
rect 6273 31457 7169 31503
rect 5618 31300 5676 31306
rect 5617 31242 5618 31300
rect 5676 31242 5975 31300
rect 5618 31234 5676 31240
rect 5677 30970 5735 30973
rect 4896 30967 5735 30970
rect 4896 30933 5689 30967
rect 5723 30933 5735 30967
rect 6273 30964 6319 31457
rect 6706 31360 6766 31366
rect 6536 31300 6706 31360
rect 6536 31254 6596 31300
rect 6706 31294 6766 31300
rect 4896 30930 5735 30933
rect 4896 29800 4936 30930
rect 5677 30927 5735 30930
rect 6272 30958 6320 30964
rect 6272 30922 6278 30958
rect 6314 30922 6320 30958
rect 6272 30916 6320 30922
rect 6273 30887 6319 30916
rect 7123 30903 7169 31457
rect 7493 31443 7539 32507
rect 8886 32510 8926 34780
rect 9446 33270 12016 33310
rect 9446 32510 9486 33270
rect 10956 32979 11186 32980
rect 10283 32978 11186 32979
rect 10283 32921 10736 32978
rect 10283 32722 10341 32921
rect 10730 32920 10736 32921
rect 10796 32921 11186 32978
rect 10796 32920 10802 32921
rect 10956 32919 11186 32921
rect 11125 32724 11186 32919
rect 10516 32540 10866 32550
rect 10516 32510 10534 32540
rect 8886 32470 9816 32510
rect 10522 32500 10534 32510
rect 10574 32510 10866 32540
rect 10574 32500 10586 32510
rect 10522 32494 10586 32500
rect 9761 32467 9816 32470
rect 9761 32455 10061 32467
rect 9761 32449 10075 32455
rect 9761 32437 10029 32449
rect 10017 32415 10029 32437
rect 10063 32415 10075 32449
rect 10017 32409 10075 32415
rect 10106 32443 10152 32455
rect 10106 32409 10112 32443
rect 10146 32440 10152 32443
rect 10146 32410 10221 32440
rect 10146 32409 10152 32410
rect 10106 32397 10152 32409
rect 10106 32340 10146 32397
rect 7656 32300 10146 32340
rect 7656 31610 7696 32300
rect 9758 32200 9816 32206
rect 9757 32140 9758 32198
rect 9816 32140 10157 32198
rect 9758 32134 9816 32140
rect 8606 31980 8666 31986
rect 7906 31979 8606 31980
rect 7879 31920 8606 31979
rect 7879 31714 7937 31920
rect 8606 31724 8666 31920
rect 7817 31610 7869 31616
rect 7656 31570 7823 31610
rect 7863 31570 7886 31610
rect 7817 31564 7869 31570
rect 7645 31443 7707 31445
rect 7493 31439 7707 31443
rect 7493 31401 7657 31439
rect 7695 31401 7707 31439
rect 7493 31397 7707 31401
rect 8207 31437 8399 31443
rect 8207 31403 8219 31437
rect 8253 31403 8399 31437
rect 8207 31397 8399 31403
rect 7645 31395 7707 31397
rect 7658 31190 7716 31196
rect 7657 31132 7658 31190
rect 7716 31132 7937 31190
rect 7658 31124 7716 31130
rect 8353 30903 8399 31397
rect 8615 31017 8676 31176
rect 8615 31011 8677 31017
rect 8615 30950 8616 31011
rect 8616 30944 8677 30950
rect 7123 30857 8399 30903
rect 5881 30660 5912 30691
rect 5917 30670 5975 30719
rect 5917 30660 6016 30670
rect 5917 30626 5975 30660
rect 5917 30620 5976 30626
rect 5917 30561 5918 30620
rect 5918 30554 5976 30560
rect 6526 30520 6586 30705
rect 6520 30460 6526 30520
rect 6586 30460 6592 30520
rect 10826 30100 10866 32510
rect 11126 32010 11186 32175
rect 11126 31944 11186 31950
rect 3826 29760 4936 29800
rect 7176 30060 10866 30100
rect 3826 28020 3866 29760
rect 4326 29310 6836 29350
rect 4326 28709 4366 29310
rect 5536 29201 5597 29207
rect 5535 29199 5536 29200
rect 4631 29141 5536 29199
rect 4631 28984 4689 29141
rect 5535 29140 5536 29141
rect 5535 29134 5597 29140
rect 5535 29004 5596 29134
rect 4323 28697 4369 28709
rect 4323 28663 4329 28697
rect 4363 28663 4369 28697
rect 4323 28651 4369 28663
rect 5057 28690 5115 28693
rect 5057 28687 5356 28690
rect 5057 28653 5069 28687
rect 5103 28653 5356 28687
rect 5057 28650 5356 28653
rect 5057 28647 5115 28650
rect 4867 28580 4925 28583
rect 4867 28577 5166 28580
rect 4867 28543 4879 28577
rect 4913 28543 5166 28577
rect 4867 28540 5166 28543
rect 4867 28537 4925 28540
rect 4631 28356 4689 28460
rect 4628 28350 4689 28356
rect 4686 28291 4689 28350
rect 4628 28284 4686 28290
rect 5126 28020 5166 28540
rect 5316 28260 5356 28650
rect 5526 28410 5586 28455
rect 5696 28410 5756 28416
rect 5526 28350 5696 28410
rect 5696 28344 5756 28350
rect 5316 28220 6286 28260
rect 3826 27980 5166 28020
rect 6246 27810 6286 28220
rect 6796 28230 6836 29310
rect 7176 28772 7216 30060
rect 7550 29280 7556 29281
rect 7406 29279 7556 29280
rect 7397 29220 7556 29279
rect 7617 29280 7623 29281
rect 7617 29220 8056 29280
rect 7397 29219 8056 29220
rect 7397 29032 7455 29219
rect 7995 29034 8056 29219
rect 7170 28760 7222 28772
rect 7170 28720 7176 28760
rect 7216 28720 7222 28760
rect 7170 28708 7222 28720
rect 7487 28740 7545 28743
rect 7487 28737 7876 28740
rect 7487 28703 7499 28737
rect 7533 28703 7876 28737
rect 7487 28700 7876 28703
rect 7487 28697 7545 28700
rect 7178 28510 7236 28516
rect 7177 28450 7178 28508
rect 7236 28450 7455 28508
rect 7178 28444 7236 28450
rect 7836 28230 7876 28700
rect 7996 28390 8056 28485
rect 8536 28430 8576 30060
rect 11976 29710 12016 33270
rect 9086 29670 12016 29710
rect 9086 29010 9126 29670
rect 9086 28970 10846 29010
rect 8870 28436 8922 28442
rect 8536 28390 8870 28430
rect 7997 28340 8056 28390
rect 8870 28378 8922 28384
rect 7990 28281 7996 28340
rect 8056 28281 8062 28340
rect 6796 28190 7876 28230
rect 9086 27810 9126 28970
rect 10436 28870 10494 28876
rect 10433 28810 10436 28869
rect 10433 28804 10494 28810
rect 10433 28614 10491 28804
rect 9290 28436 9342 28442
rect 9342 28390 10066 28430
rect 9290 28378 9342 28384
rect 10026 28339 10066 28390
rect 10806 28339 10846 28970
rect 11196 28870 11256 28876
rect 11196 28624 11256 28810
rect 10023 28327 10069 28339
rect 10023 28293 10029 28327
rect 10063 28293 10069 28327
rect 10023 28281 10069 28293
rect 10803 28327 10849 28339
rect 10803 28293 10809 28327
rect 10843 28293 10849 28327
rect 10803 28281 10849 28293
rect 10720 28214 23686 28220
rect 10720 28166 10732 28214
rect 10780 28166 23686 28214
rect 10720 28160 23686 28166
rect 23746 28160 23752 28220
rect 10048 28090 10106 28096
rect 10047 28032 10048 28090
rect 10106 28032 10399 28090
rect 10048 28024 10106 28030
rect 11196 27950 11256 28075
rect 11196 27884 11256 27890
rect 6246 27770 9126 27810
rect 3396 27040 16356 27100
rect 16416 27040 16422 27100
rect 2756 26250 15296 26310
rect 15356 26250 15362 26310
<< via1 >>
rect 6298 35220 6356 35280
rect 6946 35310 7006 35370
rect 4778 34350 4836 34410
rect 6956 34360 7016 34420
rect 4788 33980 4846 34040
rect 4700 31894 4752 31946
rect 6726 34110 6785 34170
rect 8476 34600 8536 34660
rect 8026 34420 8086 34480
rect 7538 33860 7596 33920
rect 8466 33660 8526 33720
rect 5138 33240 5196 33300
rect 6726 33270 6786 33330
rect 5908 32410 5966 32470
rect 5120 31894 5172 31946
rect 6726 32370 6785 32430
rect 5118 31510 5176 31570
rect 6726 31590 6786 31650
rect 5618 31240 5676 31300
rect 6706 31300 6766 31360
rect 10736 32920 10796 32978
rect 9758 32140 9816 32200
rect 8606 31920 8666 31980
rect 7658 31130 7716 31190
rect 8616 30950 8677 31011
rect 5918 30560 5976 30620
rect 6526 30460 6586 30520
rect 11126 31950 11186 32010
rect 5536 29140 5597 29201
rect 4628 28290 4686 28350
rect 5696 28350 5756 28410
rect 7556 29220 7617 29281
rect 7178 28450 7236 28510
rect 8870 28384 8922 28436
rect 7996 28281 8056 28340
rect 10436 28810 10494 28870
rect 9290 28384 9342 28436
rect 11196 28810 11256 28870
rect 23686 28160 23746 28220
rect 10048 28030 10106 28090
rect 11196 27890 11256 27950
rect 16356 27040 16416 27100
rect 15296 26250 15356 26310
<< metal2 >>
rect 6818 35370 6874 35377
rect 6816 35368 6946 35370
rect 6816 35312 6818 35368
rect 6874 35312 6946 35368
rect 6816 35310 6946 35312
rect 7006 35310 7012 35370
rect 6818 35303 6874 35310
rect 6158 35280 6214 35287
rect 6156 35278 6298 35280
rect 6156 35222 6158 35278
rect 6214 35222 6298 35278
rect 6156 35220 6298 35222
rect 6356 35220 6362 35280
rect 6158 35213 6214 35220
rect 8308 34660 8364 34667
rect 8306 34658 8476 34660
rect 8306 34602 8308 34658
rect 8364 34602 8476 34658
rect 8306 34600 8476 34602
rect 8536 34600 8542 34660
rect 8308 34593 8364 34600
rect 8208 34480 8264 34487
rect 8020 34420 8026 34480
rect 8086 34478 8264 34480
rect 8086 34422 8208 34478
rect 8086 34420 8264 34422
rect 3598 34410 3654 34417
rect 3596 34408 4778 34410
rect 3596 34352 3598 34408
rect 3654 34352 4778 34408
rect 3596 34350 4778 34352
rect 4836 34350 4842 34410
rect 6316 34360 6956 34420
rect 7016 34360 7022 34420
rect 8208 34413 8264 34420
rect 3598 34343 3654 34350
rect 3598 34040 3654 34047
rect 3596 34038 4788 34040
rect 3596 33982 3598 34038
rect 3654 33982 4018 34038
rect 4074 33982 4788 34038
rect 3596 33980 4788 33982
rect 4846 33980 4852 34040
rect 3598 33973 3654 33980
rect 6316 33330 6376 34360
rect 6918 34170 6974 34177
rect 6720 34110 6726 34170
rect 6785 34168 6976 34170
rect 6785 34112 6918 34168
rect 6974 34112 6976 34168
rect 6785 34110 6976 34112
rect 6918 34103 6974 34110
rect 7146 33860 7538 33920
rect 7596 33860 7602 33920
rect 7146 33720 7206 33860
rect 7146 33660 8466 33720
rect 8526 33660 8532 33720
rect 3818 33300 3874 33307
rect 3816 33298 5138 33300
rect 3816 33242 3818 33298
rect 3874 33242 5138 33298
rect 3816 33240 5138 33242
rect 5196 33240 5202 33300
rect 6316 33270 6726 33330
rect 6786 33270 6792 33330
rect 3818 33233 3874 33240
rect 4206 32860 4266 33240
rect 6316 32860 6376 33270
rect 7146 32860 7206 33660
rect 10736 33158 10796 33160
rect 10729 33102 10738 33158
rect 10794 33102 10803 33158
rect 10736 32978 10796 33102
rect 10736 32914 10796 32920
rect 4206 32800 7206 32860
rect 4206 31570 4266 32800
rect 5758 32470 5814 32477
rect 5756 32468 5908 32470
rect 5756 32412 5758 32468
rect 5814 32412 5908 32468
rect 5756 32410 5908 32412
rect 5966 32410 5972 32470
rect 5758 32403 5814 32410
rect 6720 32370 6726 32430
rect 6785 32428 6996 32430
rect 6785 32372 6938 32428
rect 6994 32372 7003 32428
rect 6785 32370 6996 32372
rect 7146 32200 7206 32800
rect 7146 32140 9758 32200
rect 9816 32140 9822 32200
rect 4694 31894 4700 31946
rect 4752 31940 4758 31946
rect 5114 31940 5120 31946
rect 4752 31900 5120 31940
rect 4752 31894 4758 31900
rect 5114 31894 5120 31900
rect 5172 31894 5178 31946
rect 7146 31650 7206 32140
rect 9446 32010 9506 32140
rect 8600 31920 8606 31980
rect 8666 31978 8846 31980
rect 8666 31922 8788 31978
rect 8844 31922 8853 31978
rect 9446 31950 11126 32010
rect 11186 31950 11192 32010
rect 8666 31920 8846 31922
rect 6720 31590 6726 31650
rect 6786 31590 7206 31650
rect 4206 31510 5118 31570
rect 5176 31510 5182 31570
rect 4206 30620 4266 31510
rect 6700 31300 6706 31360
rect 6766 31358 6936 31360
rect 6766 31302 6878 31358
rect 6934 31302 6943 31358
rect 6766 31300 6936 31302
rect 5386 31298 5618 31300
rect 5379 31242 5388 31298
rect 5444 31242 5618 31298
rect 5386 31240 5618 31242
rect 5676 31240 5682 31300
rect 7146 31190 7206 31590
rect 7146 31130 7658 31190
rect 7716 31130 7722 31190
rect 7486 31010 7546 31130
rect 8610 31010 8616 31011
rect 7486 30950 8616 31010
rect 8677 30950 8683 31011
rect 4206 30560 5918 30620
rect 5976 30560 5982 30620
rect 4206 28350 4266 30560
rect 5746 30350 5806 30560
rect 6526 30520 6586 30526
rect 6526 30350 6586 30460
rect 5746 30290 6586 30350
rect 7558 29480 7614 29487
rect 7556 29478 7616 29480
rect 7556 29422 7558 29478
rect 7614 29422 7616 29478
rect 7556 29287 7616 29422
rect 7556 29281 7617 29287
rect 7556 29214 7617 29220
rect 5530 29140 5536 29201
rect 5597 29200 5603 29201
rect 5597 29198 5806 29200
rect 5597 29142 5748 29198
rect 5804 29142 5813 29198
rect 5597 29140 5806 29142
rect 10430 28810 10436 28870
rect 10494 28868 11196 28870
rect 10494 28812 10978 28868
rect 11034 28812 11196 28868
rect 10494 28810 11196 28812
rect 11256 28810 11262 28870
rect 6226 28450 7178 28510
rect 7236 28450 7242 28510
rect 6226 28410 6286 28450
rect 5690 28350 5696 28410
rect 5756 28350 6286 28410
rect 8864 28384 8870 28436
rect 8922 28430 8928 28436
rect 9284 28430 9290 28436
rect 8922 28390 9290 28430
rect 8922 28384 8928 28390
rect 9284 28384 9290 28390
rect 9342 28384 9348 28436
rect 4206 28290 4628 28350
rect 4686 28290 4692 28350
rect 4206 27900 4266 28290
rect 6226 28090 6286 28350
rect 7996 28340 8056 28346
rect 7996 28090 8056 28281
rect 23686 28220 23746 28226
rect 6226 28030 10048 28090
rect 10106 28030 10112 28090
rect 6226 27900 6286 28030
rect 4206 27840 6286 27900
rect 9906 27790 9966 28030
rect 10966 27890 11196 27950
rect 11256 27890 11262 27950
rect 10966 27790 11026 27890
rect 9906 27730 11026 27790
rect 16356 27100 16416 27106
rect 15296 26310 15356 26316
rect 15296 14778 15356 26250
rect 16356 15748 16416 27040
rect 23686 16718 23746 28160
rect 23686 16662 23688 16718
rect 23744 16662 23746 16718
rect 23686 16660 23746 16662
rect 23688 16653 23744 16660
rect 16356 15692 16358 15748
rect 16414 15692 16416 15748
rect 16356 15690 16416 15692
rect 16358 15683 16414 15690
rect 15296 14722 15298 14778
rect 15354 14722 15356 14778
rect 15296 14720 15356 14722
rect 15298 14713 15354 14720
<< via2 >>
rect 6818 35312 6874 35368
rect 6158 35222 6214 35278
rect 8308 34602 8364 34658
rect 8208 34422 8264 34478
rect 3598 34352 3654 34408
rect 3598 33982 3654 34038
rect 4018 33982 4074 34038
rect 6918 34112 6974 34168
rect 3818 33242 3874 33298
rect 10738 33102 10794 33158
rect 5758 32412 5814 32468
rect 6938 32372 6994 32428
rect 8788 31922 8844 31978
rect 6878 31302 6934 31358
rect 5388 31242 5444 31298
rect 7558 29422 7614 29478
rect 5748 29142 5804 29198
rect 10978 28812 11034 28868
rect 23688 16662 23744 16718
rect 16358 15692 16414 15748
rect 15298 14722 15354 14778
<< metal3 >>
rect 6136 35820 7356 35880
rect 6136 35550 6196 35820
rect 5856 35490 6576 35550
rect 5856 35280 5916 35490
rect 6516 35370 6576 35490
rect 6813 35370 6879 35373
rect 6516 35368 6879 35370
rect 6516 35312 6818 35368
rect 6874 35312 6879 35368
rect 6516 35310 6879 35312
rect 6813 35307 6879 35310
rect 6153 35280 6219 35283
rect 4016 35278 6219 35280
rect 4016 35222 6158 35278
rect 6214 35222 6219 35278
rect 4016 35220 6219 35222
rect 3593 34410 3659 34413
rect 1916 34408 3659 34410
rect 1916 34352 3598 34408
rect 3654 34352 3659 34408
rect 1916 34350 3659 34352
rect 0 33810 6 34210
rect 406 34040 412 34210
rect 1168 34040 1174 34042
rect 406 33980 1174 34040
rect 406 33810 412 33980
rect 1168 33978 1174 33980
rect 1238 33978 1244 34042
rect 1916 33630 1976 34350
rect 3593 34347 3659 34350
rect 2224 34042 2288 34048
rect 4016 34043 4076 35220
rect 6153 35217 6219 35220
rect 7296 35010 7356 35820
rect 7296 34950 8196 35010
rect 7296 34440 7356 34950
rect 8136 34900 8196 34950
rect 8136 34840 8726 34900
rect 8136 34660 8196 34840
rect 8303 34660 8369 34663
rect 8136 34658 8369 34660
rect 8136 34602 8308 34658
rect 8364 34602 8369 34658
rect 8136 34600 8369 34602
rect 8303 34597 8369 34600
rect 7046 34380 7356 34440
rect 8203 34480 8269 34483
rect 8666 34480 8726 34840
rect 8203 34478 8726 34480
rect 8203 34422 8208 34478
rect 8264 34422 8726 34478
rect 8203 34420 8726 34422
rect 8203 34417 8269 34420
rect 6913 34170 6979 34173
rect 7046 34170 7106 34380
rect 6913 34168 7106 34170
rect 6913 34112 6918 34168
rect 6974 34112 7106 34168
rect 6913 34110 7106 34112
rect 6913 34107 6979 34110
rect 3593 34040 3659 34043
rect 2288 34038 3659 34040
rect 2288 33982 3598 34038
rect 3654 33982 3659 34038
rect 2288 33980 3659 33982
rect 2224 33972 2288 33978
rect 3156 33700 3216 33980
rect 3593 33977 3659 33980
rect 4013 34038 4079 34043
rect 4013 33982 4018 34038
rect 4074 33982 4079 34038
rect 4013 33977 4079 33982
rect 3156 33640 4646 33700
rect 1916 33570 2616 33630
rect 600 33070 606 33470
rect 1006 33300 1012 33470
rect 2556 33300 2616 33570
rect 3813 33300 3879 33303
rect 1006 33298 3879 33300
rect 1006 33242 3818 33298
rect 3874 33242 3879 33298
rect 1006 33240 3879 33242
rect 1006 33070 1012 33240
rect 3813 33237 3879 33240
rect 4586 32470 4646 33640
rect 8356 33370 10796 33430
rect 8356 32640 8416 33370
rect 10736 33163 10796 33370
rect 10733 33158 10799 33163
rect 10733 33102 10738 33158
rect 10794 33102 10799 33158
rect 10733 33097 10799 33102
rect 5596 32580 8846 32640
rect 5596 32470 5656 32580
rect 5753 32470 5819 32473
rect 4586 32468 5819 32470
rect 4586 32412 5758 32468
rect 5814 32412 5819 32468
rect 6936 32433 6996 32580
rect 4586 32410 5819 32412
rect 5386 31480 5446 32410
rect 5753 32407 5819 32410
rect 6933 32428 6999 32433
rect 6933 32372 6938 32428
rect 6994 32372 6999 32428
rect 6933 32367 6999 32372
rect 8786 31983 8846 32580
rect 8783 31978 8849 31983
rect 8783 31922 8788 31978
rect 8844 31922 8849 31978
rect 8783 31917 8849 31922
rect 5986 31510 6936 31570
rect 5986 31480 6046 31510
rect 5116 31420 6046 31480
rect 5116 29830 5176 31420
rect 5386 31303 5446 31420
rect 6876 31363 6936 31510
rect 6873 31358 6939 31363
rect 5383 31298 5449 31303
rect 5383 31242 5388 31298
rect 5444 31242 5449 31298
rect 6873 31302 6878 31358
rect 6934 31302 6939 31358
rect 6873 31297 6939 31302
rect 5383 31237 5449 31242
rect 6196 30220 8696 30280
rect 6196 29830 6256 30220
rect 5116 29770 6566 29830
rect 5116 29440 5176 29770
rect 6506 29480 6566 29770
rect 7553 29480 7619 29483
rect 6506 29478 7619 29480
rect 5116 29380 5806 29440
rect 6506 29422 7558 29478
rect 7614 29422 7619 29478
rect 6506 29420 7619 29422
rect 7553 29417 7619 29420
rect 5746 29203 5806 29380
rect 8636 29350 8696 30220
rect 8636 29290 11036 29350
rect 5743 29198 5809 29203
rect 5743 29142 5748 29198
rect 5804 29142 5809 29198
rect 5743 29137 5809 29142
rect 10976 28873 11036 29290
rect 10973 28868 11039 28873
rect 10973 28812 10978 28868
rect 11034 28812 11039 28868
rect 10973 28807 11039 28812
rect 23683 16720 23749 16723
rect 23683 16718 29586 16720
rect 23683 16662 23688 16718
rect 23744 16662 29586 16718
rect 23683 16660 29586 16662
rect 23683 16657 23749 16660
rect 16353 15750 16419 15753
rect 16353 15748 25556 15750
rect 16353 15692 16358 15748
rect 16414 15692 25556 15748
rect 16353 15690 25556 15692
rect 16353 15687 16419 15690
rect 15293 14780 15359 14783
rect 15293 14778 21786 14780
rect 15293 14722 15298 14778
rect 15354 14722 21786 14778
rect 15293 14720 21786 14722
rect 15293 14717 15359 14720
rect 21726 720 21786 14720
rect 21726 660 22056 720
rect 21996 340 22056 660
rect 25496 390 25556 15690
rect 29526 800 29586 16660
rect 29526 740 30286 800
rect 21996 280 22556 340
rect 25496 330 26426 390
rect 22496 206 22556 280
rect 22436 200 22616 206
rect 26366 196 26426 330
rect 30226 196 30286 740
rect 22436 14 22616 20
rect 26306 190 26486 196
rect 26306 4 26486 10
rect 30166 190 30346 196
rect 30166 4 30346 10
<< via3 >>
rect 6 33810 406 34210
rect 1174 33978 1238 34042
rect 2224 33978 2288 34042
rect 606 33070 1006 33470
rect 22436 20 22616 200
rect 26306 10 26486 190
rect 30166 10 30346 190
<< metal4 >>
rect 5940 44952 6000 45152
rect 6492 44952 6552 45152
rect 7044 44952 7104 45152
rect 7596 44952 7656 45152
rect 8148 44952 8208 45152
rect 8700 44952 8760 45152
rect 9252 44952 9312 45152
rect 9804 44952 9864 45152
rect 10356 44952 10416 45152
rect 10908 44952 10968 45152
rect 11460 44952 11520 45152
rect 12012 44952 12072 45152
rect 12564 44952 12624 45152
rect 13116 44952 13176 45152
rect 13668 44952 13728 45152
rect 14220 44952 14280 45152
rect 14772 44952 14832 45152
rect 15324 44952 15384 45152
rect 15876 44952 15936 45152
rect 16428 44952 16488 45152
rect 16980 44952 17040 45152
rect 17532 44952 17592 45152
rect 18084 44952 18144 45152
rect 18636 44952 18696 45152
rect 19188 44952 19248 45152
rect 19740 44952 19800 45152
rect 20292 44952 20352 45152
rect 20844 44952 20904 45152
rect 21396 44952 21456 45152
rect 21948 44952 22008 45152
rect 22500 44952 22560 45152
rect 23052 44952 23112 45152
rect 23604 44952 23664 45152
rect 24156 44952 24216 45152
rect 24708 44952 24768 45152
rect 25260 44952 25320 45152
rect 25812 44952 25872 45152
rect 26364 44952 26424 45152
rect 26916 44952 26976 45152
rect 27468 44952 27528 45152
rect 28020 44952 28080 45152
rect 28572 44952 28632 45152
rect 29124 44952 29184 45152
rect 6 34211 406 44152
rect 5 34210 407 34211
rect 5 33810 6 34210
rect 406 33810 407 34210
rect 5 33809 407 33810
rect 6 1000 406 33809
rect 606 33471 1006 44152
rect 1173 34042 1239 34043
rect 1173 33978 1174 34042
rect 1238 34040 1239 34042
rect 2223 34042 2289 34043
rect 2223 34040 2224 34042
rect 1238 33980 2224 34040
rect 1238 33978 1239 33980
rect 1173 33977 1239 33978
rect 2223 33978 2224 33980
rect 2288 33978 2289 34042
rect 2223 33977 2289 33978
rect 605 33470 1007 33471
rect 605 33070 606 33470
rect 1006 33070 1007 33470
rect 605 33069 1007 33070
rect 606 1000 1006 33069
rect 22435 200 22617 201
rect 3120 0 3300 200
rect 6984 0 7164 200
rect 10848 0 11028 200
rect 14712 0 14892 200
rect 18576 0 18756 200
rect 22435 20 22436 200
rect 22616 20 22620 200
rect 22435 19 22620 20
rect 22440 0 22620 19
rect 26304 191 26484 200
rect 30168 191 30348 200
rect 26304 190 26487 191
rect 26304 10 26306 190
rect 26486 10 26487 190
rect 26304 9 26487 10
rect 30165 190 30348 191
rect 30165 10 30166 190
rect 30346 10 30348 190
rect 30165 9 30348 10
rect 26304 0 26484 9
rect 30168 0 30348 9
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8 ~/sky130_skel
timestamp 1731027661
transform 1 0 5514 0 1 28458
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 /edatools/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731131477
transform 1 0 4476 0 1 28450
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4 /edatools/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731131477
transform 1 0 7334 0 1 28498
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1731027661
transform 1 0 7984 0 1 28488
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_1
timestamp 1731131477
transform 1 0 10186 0 1 28080
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1731027661
transform 1 0 11184 0 1 28078
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1731131477
transform 1 0 5854 0 1 30708
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1731027661
transform 1 0 6514 0 1 30708
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1 /edatools/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731131477
transform 1 0 7816 0 1 31180
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1731027661
transform 1 0 8594 0 1 31178
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1731131477
transform 1 0 5846 0 1 31680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1731027661
transform 1 0 6544 0 1 31688
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0 /edatools/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731131477
transform 1 0 9944 0 1 32188
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1731027661
transform 1 0 11114 0 1 32178
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1731131477
transform 1 0 6056 0 1 33450
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1731027661
transform 1 0 6714 0 1 33448
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1731131477
transform 1 0 7666 0 1 33910
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1731027661
transform 1 0 8456 0 1 33850
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1731131477
transform 1 0 6146 0 1 34510
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1731027661
transform 1 0 6934 0 1 34508
box -38 -48 130 592
<< labels >>
rlabel metal4 s 28572 44952 28632 45152 6 clk
port 0 nsew default input
rlabel metal4 s 29124 44952 29184 45152 6 ena
port 1 nsew default input
rlabel metal4 s 28020 44952 28080 45152 6 rst_n
port 2 nsew default input
rlabel metal4 s 30168 0 30348 200 6 ua[0]
port 3 nsew default bidirectional
rlabel metal4 s 26304 0 26484 200 6 ua[1]
port 4 nsew default bidirectional
rlabel metal4 s 22440 0 22620 200 6 ua[2]
port 5 nsew default bidirectional
rlabel metal4 s 18576 0 18756 200 6 ua[3]
port 6 nsew default bidirectional
rlabel metal4 s 14712 0 14892 200 6 ua[4]
port 7 nsew default bidirectional
rlabel metal4 s 10848 0 11028 200 6 ua[5]
port 8 nsew default bidirectional
rlabel metal4 s 6984 0 7164 200 6 ua[6]
port 9 nsew default bidirectional
rlabel metal4 s 3120 0 3300 200 6 ua[7]
port 10 nsew default bidirectional
rlabel metal4 s 27468 44952 27528 45152 6 ui_in[0]
port 11 nsew default input
rlabel metal4 s 26916 44952 26976 45152 6 ui_in[1]
port 12 nsew default input
rlabel metal4 s 26364 44952 26424 45152 6 ui_in[2]
port 13 nsew default input
rlabel metal4 s 25812 44952 25872 45152 6 ui_in[3]
port 14 nsew default input
rlabel metal4 s 25260 44952 25320 45152 6 ui_in[4]
port 15 nsew default input
rlabel metal4 s 24708 44952 24768 45152 6 ui_in[5]
port 16 nsew default input
rlabel metal4 s 24156 44952 24216 45152 6 ui_in[6]
port 17 nsew default input
rlabel metal4 s 23604 44952 23664 45152 6 ui_in[7]
port 18 nsew default input
rlabel metal4 s 23052 44952 23112 45152 6 uio_in[0]
port 19 nsew default input
rlabel metal4 s 22500 44952 22560 45152 6 uio_in[1]
port 20 nsew default input
rlabel metal4 s 21948 44952 22008 45152 6 uio_in[2]
port 21 nsew default input
rlabel metal4 s 21396 44952 21456 45152 6 uio_in[3]
port 22 nsew default input
rlabel metal4 s 20844 44952 20904 45152 6 uio_in[4]
port 23 nsew default input
rlabel metal4 s 20292 44952 20352 45152 6 uio_in[5]
port 24 nsew default input
rlabel metal4 s 19740 44952 19800 45152 6 uio_in[6]
port 25 nsew default input
rlabel metal4 s 19188 44952 19248 45152 6 uio_in[7]
port 26 nsew default input
rlabel metal4 s 9804 44952 9864 45152 6 uio_oe[0]
port 27 nsew default tristate
rlabel metal4 s 9252 44952 9312 45152 6 uio_oe[1]
port 28 nsew default tristate
rlabel metal4 s 8700 44952 8760 45152 6 uio_oe[2]
port 29 nsew default tristate
rlabel metal4 s 8148 44952 8208 45152 6 uio_oe[3]
port 30 nsew default tristate
rlabel metal4 s 7596 44952 7656 45152 6 uio_oe[4]
port 31 nsew default tristate
rlabel metal4 s 7044 44952 7104 45152 6 uio_oe[5]
port 32 nsew default tristate
rlabel metal4 s 6492 44952 6552 45152 6 uio_oe[6]
port 33 nsew default tristate
rlabel metal4 s 5940 44952 6000 45152 6 uio_oe[7]
port 34 nsew default tristate
rlabel metal4 s 14220 44952 14280 45152 6 uio_out[0]
port 35 nsew default tristate
rlabel metal4 s 13668 44952 13728 45152 6 uio_out[1]
port 36 nsew default tristate
rlabel metal4 s 13116 44952 13176 45152 6 uio_out[2]
port 37 nsew default tristate
rlabel metal4 s 12564 44952 12624 45152 6 uio_out[3]
port 38 nsew default tristate
rlabel metal4 s 12012 44952 12072 45152 6 uio_out[4]
port 39 nsew default tristate
rlabel metal4 s 11460 44952 11520 45152 6 uio_out[5]
port 40 nsew default tristate
rlabel metal4 s 10908 44952 10968 45152 6 uio_out[6]
port 41 nsew default tristate
rlabel metal4 s 10356 44952 10416 45152 6 uio_out[7]
port 42 nsew default tristate
rlabel metal4 s 18636 44952 18696 45152 6 uo_out[0]
port 43 nsew default tristate
rlabel metal4 s 18084 44952 18144 45152 6 uo_out[1]
port 44 nsew default tristate
rlabel metal4 s 17532 44952 17592 45152 6 uo_out[2]
port 45 nsew default tristate
rlabel metal4 s 16980 44952 17040 45152 6 uo_out[3]
port 46 nsew default tristate
rlabel metal4 s 16428 44952 16488 45152 6 uo_out[4]
port 47 nsew default tristate
rlabel metal4 s 15876 44952 15936 45152 6 uo_out[5]
port 48 nsew default tristate
rlabel metal4 s 15324 44952 15384 45152 6 uo_out[6]
port 49 nsew default tristate
rlabel metal4 s 14772 44952 14832 45152 6 uo_out[7]
port 50 nsew default tristate
flabel metal4 6 1000 406 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 606 1000 1006 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< end >>
