magic
tech sky130A
magscale 1 2
timestamp 1731266928
<< nwell >>
rect 6333 35090 6910 35092
rect 6333 34771 7258 35090
rect 6906 34769 7258 34771
rect 7853 34432 8430 34492
rect 7853 34171 8780 34432
rect 8426 34111 8780 34171
rect 6243 34030 6730 34032
rect 6243 33711 7038 34030
rect 6726 33709 7038 33711
rect 10499 32760 11080 32770
rect 10499 32449 11438 32760
rect 11066 32439 11438 32449
rect 6526 32262 6868 32270
rect 6033 31949 6868 32262
rect 6033 31941 6550 31949
rect 8003 31760 8580 31762
rect 8003 31441 8918 31760
rect 8576 31439 8918 31441
rect 6041 30969 6838 31290
rect 7521 29070 8010 29080
rect 5506 29032 5838 29040
rect 4847 28719 5838 29032
rect 7521 28759 8308 29070
rect 7976 28749 8308 28759
rect 4847 28711 5510 28719
rect 10557 28660 11160 28662
rect 10557 28341 11508 28660
rect 11156 28339 11508 28341
<< locali >>
rect 6200 34767 6432 34770
rect 6200 34733 6203 34767
rect 6237 34733 6432 34767
rect 6200 34730 6432 34733
rect 6504 34737 6823 34743
rect 6504 34703 6783 34737
rect 6817 34703 6823 34737
rect 6504 34697 6823 34703
rect 7730 34617 7860 34620
rect 7730 34583 7813 34617
rect 7847 34583 7860 34617
rect 7730 34580 7860 34583
rect 7730 34350 7770 34580
rect 7730 34310 7940 34350
rect 8090 34167 8359 34169
rect 8090 34133 8323 34167
rect 8357 34133 8359 34167
rect 8090 34131 8359 34133
rect 6090 33707 6342 33710
rect 6090 33673 6093 33707
rect 6127 33673 6342 33707
rect 6090 33670 6342 33673
rect 6414 33677 6713 33683
rect 6414 33643 6673 33677
rect 6707 33643 6713 33677
rect 6414 33637 6713 33643
rect 10731 32550 10765 32563
rect 10731 32540 10780 32550
rect 10768 32500 10780 32540
rect 10760 32490 10780 32500
rect 10223 32449 10272 32486
rect 10257 32415 10272 32449
rect 10223 32406 10272 32415
rect 10340 32409 10407 32443
rect 5870 31937 6132 31940
rect 5870 31903 5873 31937
rect 5907 31903 6132 31937
rect 5870 31900 6132 31903
rect 6204 31877 6513 31903
rect 6204 31857 6473 31877
rect 6467 31843 6473 31857
rect 6507 31843 6513 31877
rect 6467 31827 6513 31843
rect 8000 31610 8030 31620
rect 8000 31570 8017 31610
rect 8000 31560 8030 31570
rect 7815 31439 8047 31445
rect 7815 31401 7851 31439
rect 7889 31401 8047 31439
rect 8140 31412 8156 31460
rect 8226 31440 8242 31445
rect 8226 31437 8460 31440
rect 8226 31403 8413 31437
rect 8447 31403 8460 31437
rect 8226 31402 8460 31403
rect 7815 31395 8047 31401
rect 8239 31400 8460 31402
rect 5880 30967 6140 30970
rect 5880 30933 5883 30967
rect 5917 30933 6140 30967
rect 6467 30958 6513 30983
rect 6467 30933 6472 30958
rect 5880 30930 6140 30933
rect 6212 30922 6472 30933
rect 6508 30922 6513 30958
rect 6212 30887 6513 30922
rect 7410 28720 7600 28760
rect 4520 28697 4717 28700
rect 4520 28663 4523 28697
rect 4557 28663 4717 28697
rect 4520 28660 4717 28663
rect 5086 28687 5300 28690
rect 5086 28653 5263 28687
rect 5297 28653 5300 28687
rect 5086 28650 5300 28653
rect 10220 28329 10400 28330
rect 10220 28327 10427 28329
rect 10220 28293 10223 28327
rect 10257 28293 10427 28327
rect 10220 28290 10427 28293
rect 10796 28327 11040 28330
rect 10796 28293 11003 28327
rect 11037 28293 11040 28327
rect 10796 28290 11040 28293
rect 10776 28214 10980 28220
rect 10776 28166 10926 28214
rect 10974 28166 10980 28214
rect 10776 28160 10980 28166
<< viali >>
rect 6203 34733 6237 34767
rect 6783 34703 6817 34737
rect 7813 34583 7847 34617
rect 7903 34133 7937 34167
rect 8323 34133 8357 34167
rect 6093 33673 6127 33707
rect 6673 33643 6707 33677
rect 10728 32500 10768 32540
rect 10223 32415 10257 32449
rect 10306 32409 10340 32443
rect 5873 31903 5907 31937
rect 6473 31843 6507 31877
rect 8017 31570 8057 31610
rect 7851 31401 7889 31439
rect 8413 31403 8447 31437
rect 5883 30933 5917 30967
rect 6472 30922 6508 30958
rect 7370 28720 7410 28760
rect 7693 28703 7727 28737
rect 4523 28663 4557 28697
rect 5263 28653 5297 28687
rect 5073 28543 5107 28577
rect 10223 28293 10257 28327
rect 11003 28293 11037 28327
rect 10926 28166 10974 28214
<< metal1 >>
rect 6777 35657 7673 35703
rect 6492 35280 6550 35286
rect 6550 35220 6553 35279
rect 6492 35214 6553 35220
rect 6495 35044 6553 35214
rect 6191 34770 6249 34773
rect 2950 34767 6249 34770
rect 2950 34733 6203 34767
rect 6237 34733 6249 34767
rect 2950 34730 6249 34733
rect 2950 26310 3010 34730
rect 6191 34727 6249 34730
rect 6777 34737 6823 35657
rect 7140 35370 7200 35376
rect 7140 35054 7200 35310
rect 6777 34703 6783 34737
rect 6817 34703 6823 34737
rect 6777 34691 6823 34703
rect 4972 34410 5030 34416
rect 4971 34351 4972 34409
rect 6403 34409 6461 34520
rect 5030 34351 6461 34409
rect 7150 34420 7210 34505
rect 7150 34354 7210 34360
rect 4972 34344 5030 34350
rect 6667 34237 7473 34283
rect 5841 34131 6371 34189
rect 4982 34040 5040 34046
rect 4981 33981 4982 34039
rect 5841 34039 5899 34131
rect 5040 33981 5899 34039
rect 6313 33984 6371 34131
rect 4982 33974 5040 33980
rect 6081 33710 6139 33713
rect 5090 33707 6139 33710
rect 5090 33673 6093 33707
rect 6127 33673 6139 33707
rect 5090 33670 6139 33673
rect 4894 31946 4946 31952
rect 3590 31900 4894 31940
rect 3590 27100 3650 31900
rect 4894 31888 4946 31894
rect 5090 30970 5130 33670
rect 6081 33667 6139 33670
rect 6667 33677 6713 34237
rect 6920 34170 6979 34176
rect 6920 33995 6979 34110
rect 7427 33733 7473 34237
rect 7627 34173 7673 35657
rect 8210 34780 9120 34820
rect 7801 34620 7859 34623
rect 8210 34620 8250 34780
rect 8670 34660 8730 34666
rect 7800 34617 8250 34620
rect 7800 34583 7813 34617
rect 7847 34583 8250 34617
rect 7800 34580 8250 34583
rect 8669 34600 8670 34660
rect 8669 34594 8730 34600
rect 7801 34577 7859 34580
rect 8220 34480 8280 34486
rect 8130 34420 8220 34480
rect 8220 34414 8280 34420
rect 8669 34396 8729 34594
rect 7627 34167 7949 34173
rect 7627 34133 7903 34167
rect 7937 34133 7949 34167
rect 7627 34127 7949 34133
rect 8317 34167 8363 34179
rect 8317 34133 8323 34167
rect 8357 34133 8363 34167
rect 7732 33920 7790 33926
rect 7731 33862 7732 33920
rect 7790 33862 7981 33920
rect 7732 33854 7790 33860
rect 8317 33733 8363 34133
rect 7427 33687 8363 33733
rect 8660 33720 8720 33847
rect 6667 33643 6673 33677
rect 6707 33643 6713 33677
rect 8660 33654 8720 33660
rect 6667 33631 6713 33643
rect 5332 33300 5390 33306
rect 5331 33241 5332 33299
rect 6313 33299 6371 33460
rect 5390 33241 6371 33299
rect 6919 33336 6979 33445
rect 6919 33330 6980 33336
rect 6919 33270 6920 33330
rect 6920 33264 6980 33270
rect 5332 33234 5390 33240
rect 6467 32507 7733 32553
rect 6102 32470 6160 32476
rect 6160 32410 6161 32469
rect 6102 32404 6161 32410
rect 6103 32214 6161 32404
rect 5314 31946 5366 31952
rect 5861 31940 5919 31943
rect 5366 31937 5919 31940
rect 5366 31903 5873 31937
rect 5907 31903 5919 31937
rect 5366 31900 5919 31903
rect 5861 31897 5919 31900
rect 5314 31888 5366 31894
rect 6467 31877 6513 32507
rect 6920 32430 6979 32436
rect 6750 32370 6920 32429
rect 6750 32235 6809 32370
rect 6920 32364 6979 32370
rect 6467 31843 6473 31877
rect 6507 31843 6513 31877
rect 6467 31831 6513 31843
rect 5312 31570 5370 31576
rect 5311 31511 5312 31569
rect 6103 31569 6161 31690
rect 6749 31650 6809 31685
rect 6920 31650 6980 31656
rect 6749 31590 6920 31650
rect 6920 31584 6980 31590
rect 5370 31511 6161 31569
rect 5312 31504 5370 31510
rect 6467 31457 7363 31503
rect 5812 31300 5870 31306
rect 5811 31242 5812 31300
rect 5870 31242 6169 31300
rect 5812 31234 5870 31240
rect 5871 30970 5929 30973
rect 5090 30967 5929 30970
rect 5090 30933 5883 30967
rect 5917 30933 5929 30967
rect 6467 30964 6513 31457
rect 6900 31360 6960 31366
rect 6730 31300 6900 31360
rect 6730 31254 6790 31300
rect 6900 31294 6960 31300
rect 5090 30930 5929 30933
rect 5090 29800 5130 30930
rect 5871 30927 5929 30930
rect 6466 30958 6514 30964
rect 6466 30922 6472 30958
rect 6508 30922 6514 30958
rect 6466 30916 6514 30922
rect 6467 30887 6513 30916
rect 7317 30903 7363 31457
rect 7687 31443 7733 32507
rect 9080 32510 9120 34780
rect 9640 33270 12210 33310
rect 9640 32510 9680 33270
rect 11150 32979 11380 32980
rect 10477 32978 11380 32979
rect 10477 32921 10930 32978
rect 10477 32722 10535 32921
rect 10924 32920 10930 32921
rect 10990 32921 11380 32978
rect 10990 32920 10996 32921
rect 11150 32919 11380 32921
rect 11319 32724 11380 32919
rect 10710 32540 11060 32550
rect 10710 32510 10728 32540
rect 9080 32470 10010 32510
rect 10716 32500 10728 32510
rect 10768 32510 11060 32540
rect 10768 32500 10780 32510
rect 10716 32494 10780 32500
rect 9955 32467 10010 32470
rect 9955 32455 10255 32467
rect 9955 32449 10269 32455
rect 9955 32437 10223 32449
rect 10211 32415 10223 32437
rect 10257 32415 10269 32449
rect 10211 32409 10269 32415
rect 10300 32443 10346 32455
rect 10300 32409 10306 32443
rect 10340 32440 10346 32443
rect 10340 32410 10415 32440
rect 10340 32409 10346 32410
rect 10300 32397 10346 32409
rect 10300 32340 10340 32397
rect 7850 32300 10340 32340
rect 7850 31610 7890 32300
rect 9952 32200 10010 32206
rect 9951 32140 9952 32198
rect 10010 32140 10351 32198
rect 9952 32134 10010 32140
rect 8800 31980 8860 31986
rect 8100 31979 8800 31980
rect 8073 31920 8800 31979
rect 8073 31714 8131 31920
rect 8800 31724 8860 31920
rect 8011 31610 8063 31616
rect 7850 31570 8017 31610
rect 8057 31570 8080 31610
rect 8011 31564 8063 31570
rect 7839 31443 7901 31445
rect 7687 31439 7901 31443
rect 7687 31401 7851 31439
rect 7889 31401 7901 31439
rect 7687 31397 7901 31401
rect 8401 31437 8593 31443
rect 8401 31403 8413 31437
rect 8447 31403 8593 31437
rect 8401 31397 8593 31403
rect 7839 31395 7901 31397
rect 7852 31190 7910 31196
rect 7851 31132 7852 31190
rect 7910 31132 8131 31190
rect 7852 31124 7910 31130
rect 8547 30903 8593 31397
rect 8809 31017 8870 31176
rect 8809 31011 8871 31017
rect 8809 30950 8810 31011
rect 8810 30944 8871 30950
rect 7317 30857 8593 30903
rect 6075 30660 6106 30691
rect 6111 30670 6169 30719
rect 6111 30660 6210 30670
rect 6111 30626 6169 30660
rect 6111 30620 6170 30626
rect 6111 30561 6112 30620
rect 6112 30554 6170 30560
rect 6720 30520 6780 30705
rect 6714 30460 6720 30520
rect 6780 30460 6786 30520
rect 11020 30100 11060 32510
rect 11320 32010 11380 32175
rect 11320 31944 11380 31950
rect 4020 29760 5130 29800
rect 7370 30060 11060 30100
rect 4020 28020 4060 29760
rect 4520 29310 7030 29350
rect 4520 28709 4560 29310
rect 5730 29201 5791 29207
rect 5729 29199 5730 29200
rect 4825 29141 5730 29199
rect 4825 28984 4883 29141
rect 5729 29140 5730 29141
rect 5729 29134 5791 29140
rect 5729 29004 5790 29134
rect 4517 28697 4563 28709
rect 4517 28663 4523 28697
rect 4557 28663 4563 28697
rect 4517 28651 4563 28663
rect 5251 28690 5309 28693
rect 5251 28687 5550 28690
rect 5251 28653 5263 28687
rect 5297 28653 5550 28687
rect 5251 28650 5550 28653
rect 5251 28647 5309 28650
rect 5061 28580 5119 28583
rect 5061 28577 5360 28580
rect 5061 28543 5073 28577
rect 5107 28543 5360 28577
rect 5061 28540 5360 28543
rect 5061 28537 5119 28540
rect 4825 28356 4883 28460
rect 4822 28350 4883 28356
rect 4880 28291 4883 28350
rect 4822 28284 4880 28290
rect 5320 28020 5360 28540
rect 5510 28260 5550 28650
rect 5720 28410 5780 28455
rect 5890 28410 5950 28416
rect 5720 28350 5890 28410
rect 5890 28344 5950 28350
rect 5510 28220 6480 28260
rect 4020 27980 5360 28020
rect 6440 27810 6480 28220
rect 6990 28230 7030 29310
rect 7370 28772 7410 30060
rect 7744 29280 7750 29281
rect 7600 29279 7750 29280
rect 7591 29220 7750 29279
rect 7811 29280 7817 29281
rect 7811 29220 8250 29280
rect 7591 29219 8250 29220
rect 7591 29032 7649 29219
rect 8189 29034 8250 29219
rect 7364 28760 7416 28772
rect 7364 28720 7370 28760
rect 7410 28720 7416 28760
rect 7364 28708 7416 28720
rect 7681 28740 7739 28743
rect 7681 28737 8070 28740
rect 7681 28703 7693 28737
rect 7727 28703 8070 28737
rect 7681 28700 8070 28703
rect 7681 28697 7739 28700
rect 7372 28510 7430 28516
rect 7371 28450 7372 28508
rect 7430 28450 7649 28508
rect 7372 28444 7430 28450
rect 8030 28230 8070 28700
rect 8190 28390 8250 28485
rect 8730 28430 8770 30060
rect 12170 29710 12210 33270
rect 9280 29670 12210 29710
rect 9280 29010 9320 29670
rect 9280 28970 11040 29010
rect 9064 28436 9116 28442
rect 8730 28390 9064 28430
rect 8191 28340 8250 28390
rect 9064 28378 9116 28384
rect 8184 28281 8190 28340
rect 8250 28281 8256 28340
rect 6990 28190 8070 28230
rect 9280 27810 9320 28970
rect 10630 28870 10688 28876
rect 10627 28810 10630 28869
rect 10627 28804 10688 28810
rect 10627 28614 10685 28804
rect 9484 28436 9536 28442
rect 9536 28390 10260 28430
rect 9484 28378 9536 28384
rect 10220 28339 10260 28390
rect 11000 28339 11040 28970
rect 11390 28870 11450 28876
rect 11390 28624 11450 28810
rect 10217 28327 10263 28339
rect 10217 28293 10223 28327
rect 10257 28293 10263 28327
rect 10217 28281 10263 28293
rect 10997 28327 11043 28339
rect 10997 28293 11003 28327
rect 11037 28293 11043 28327
rect 10997 28281 11043 28293
rect 10914 28214 23880 28220
rect 10914 28166 10926 28214
rect 10974 28166 23880 28214
rect 10914 28160 23880 28166
rect 23940 28160 23946 28220
rect 10242 28090 10300 28096
rect 10241 28032 10242 28090
rect 10300 28032 10593 28090
rect 10242 28024 10300 28030
rect 11390 27950 11450 28075
rect 11390 27884 11450 27890
rect 6440 27770 9320 27810
rect 3590 27040 16550 27100
rect 16610 27040 16616 27100
rect 2950 26250 15490 26310
rect 15550 26250 15556 26310
<< via1 >>
rect 6492 35220 6550 35280
rect 7140 35310 7200 35370
rect 4972 34350 5030 34410
rect 7150 34360 7210 34420
rect 4982 33980 5040 34040
rect 4894 31894 4946 31946
rect 6920 34110 6979 34170
rect 8670 34600 8730 34660
rect 8220 34420 8280 34480
rect 7732 33860 7790 33920
rect 8660 33660 8720 33720
rect 5332 33240 5390 33300
rect 6920 33270 6980 33330
rect 6102 32410 6160 32470
rect 5314 31894 5366 31946
rect 6920 32370 6979 32430
rect 5312 31510 5370 31570
rect 6920 31590 6980 31650
rect 5812 31240 5870 31300
rect 6900 31300 6960 31360
rect 10930 32920 10990 32978
rect 9952 32140 10010 32200
rect 8800 31920 8860 31980
rect 7852 31130 7910 31190
rect 8810 30950 8871 31011
rect 6112 30560 6170 30620
rect 6720 30460 6780 30520
rect 11320 31950 11380 32010
rect 5730 29140 5791 29201
rect 4822 28290 4880 28350
rect 5890 28350 5950 28410
rect 7750 29220 7811 29281
rect 7372 28450 7430 28510
rect 9064 28384 9116 28436
rect 8190 28281 8250 28340
rect 10630 28810 10688 28870
rect 9484 28384 9536 28436
rect 11390 28810 11450 28870
rect 23880 28160 23940 28220
rect 10242 28030 10300 28090
rect 11390 27890 11450 27950
rect 16550 27040 16610 27100
rect 15490 26250 15550 26310
<< metal2 >>
rect 7012 35370 7068 35377
rect 7010 35368 7140 35370
rect 7010 35312 7012 35368
rect 7068 35312 7140 35368
rect 7010 35310 7140 35312
rect 7200 35310 7206 35370
rect 7012 35303 7068 35310
rect 6352 35280 6408 35287
rect 6350 35278 6492 35280
rect 6350 35222 6352 35278
rect 6408 35222 6492 35278
rect 6350 35220 6492 35222
rect 6550 35220 6556 35280
rect 6352 35213 6408 35220
rect 8502 34660 8558 34667
rect 8500 34658 8670 34660
rect 8500 34602 8502 34658
rect 8558 34602 8670 34658
rect 8500 34600 8670 34602
rect 8730 34600 8736 34660
rect 8502 34593 8558 34600
rect 8402 34480 8458 34487
rect 8214 34420 8220 34480
rect 8280 34478 8458 34480
rect 8280 34422 8402 34478
rect 8280 34420 8458 34422
rect 3792 34410 3848 34417
rect 3790 34408 4972 34410
rect 3790 34352 3792 34408
rect 3848 34352 4972 34408
rect 3790 34350 4972 34352
rect 5030 34350 5036 34410
rect 6510 34360 7150 34420
rect 7210 34360 7216 34420
rect 8402 34413 8458 34420
rect 3792 34343 3848 34350
rect 3792 34040 3848 34047
rect 3790 34038 4982 34040
rect 3790 33982 3792 34038
rect 3848 33982 4212 34038
rect 4268 33982 4982 34038
rect 3790 33980 4982 33982
rect 5040 33980 5046 34040
rect 3792 33973 3848 33980
rect 6510 33330 6570 34360
rect 7112 34170 7168 34177
rect 6914 34110 6920 34170
rect 6979 34168 7170 34170
rect 6979 34112 7112 34168
rect 7168 34112 7170 34168
rect 6979 34110 7170 34112
rect 7112 34103 7168 34110
rect 7340 33860 7732 33920
rect 7790 33860 7796 33920
rect 7340 33720 7400 33860
rect 7340 33660 8660 33720
rect 8720 33660 8726 33720
rect 4012 33300 4068 33307
rect 4010 33298 5332 33300
rect 4010 33242 4012 33298
rect 4068 33242 5332 33298
rect 4010 33240 5332 33242
rect 5390 33240 5396 33300
rect 6510 33270 6920 33330
rect 6980 33270 6986 33330
rect 4012 33233 4068 33240
rect 4400 32860 4460 33240
rect 6510 32860 6570 33270
rect 7340 32860 7400 33660
rect 10930 33158 10990 33160
rect 10923 33102 10932 33158
rect 10988 33102 10997 33158
rect 10930 32978 10990 33102
rect 10930 32914 10990 32920
rect 4400 32800 7400 32860
rect 4400 31570 4460 32800
rect 5952 32470 6008 32477
rect 5950 32468 6102 32470
rect 5950 32412 5952 32468
rect 6008 32412 6102 32468
rect 5950 32410 6102 32412
rect 6160 32410 6166 32470
rect 5952 32403 6008 32410
rect 6914 32370 6920 32430
rect 6979 32428 7190 32430
rect 6979 32372 7132 32428
rect 7188 32372 7197 32428
rect 6979 32370 7190 32372
rect 7340 32200 7400 32800
rect 7340 32140 9952 32200
rect 10010 32140 10016 32200
rect 4888 31894 4894 31946
rect 4946 31940 4952 31946
rect 5308 31940 5314 31946
rect 4946 31900 5314 31940
rect 4946 31894 4952 31900
rect 5308 31894 5314 31900
rect 5366 31894 5372 31946
rect 7340 31650 7400 32140
rect 9640 32010 9700 32140
rect 8794 31920 8800 31980
rect 8860 31978 9040 31980
rect 8860 31922 8982 31978
rect 9038 31922 9047 31978
rect 9640 31950 11320 32010
rect 11380 31950 11386 32010
rect 8860 31920 9040 31922
rect 6914 31590 6920 31650
rect 6980 31590 7400 31650
rect 4400 31510 5312 31570
rect 5370 31510 5376 31570
rect 4400 30620 4460 31510
rect 6894 31300 6900 31360
rect 6960 31358 7130 31360
rect 6960 31302 7072 31358
rect 7128 31302 7137 31358
rect 6960 31300 7130 31302
rect 5580 31298 5812 31300
rect 5573 31242 5582 31298
rect 5638 31242 5812 31298
rect 5580 31240 5812 31242
rect 5870 31240 5876 31300
rect 7340 31190 7400 31590
rect 7340 31130 7852 31190
rect 7910 31130 7916 31190
rect 7680 31010 7740 31130
rect 8804 31010 8810 31011
rect 7680 30950 8810 31010
rect 8871 30950 8877 31011
rect 4400 30560 6112 30620
rect 6170 30560 6176 30620
rect 4400 28350 4460 30560
rect 5940 30350 6000 30560
rect 6720 30520 6780 30526
rect 6720 30350 6780 30460
rect 5940 30290 6780 30350
rect 7752 29480 7808 29487
rect 7750 29478 7810 29480
rect 7750 29422 7752 29478
rect 7808 29422 7810 29478
rect 7750 29287 7810 29422
rect 7750 29281 7811 29287
rect 7750 29214 7811 29220
rect 5724 29140 5730 29201
rect 5791 29200 5797 29201
rect 5791 29198 6000 29200
rect 5791 29142 5942 29198
rect 5998 29142 6007 29198
rect 5791 29140 6000 29142
rect 10624 28810 10630 28870
rect 10688 28868 11390 28870
rect 10688 28812 11172 28868
rect 11228 28812 11390 28868
rect 10688 28810 11390 28812
rect 11450 28810 11456 28870
rect 6420 28450 7372 28510
rect 7430 28450 7436 28510
rect 6420 28410 6480 28450
rect 5884 28350 5890 28410
rect 5950 28350 6480 28410
rect 9058 28384 9064 28436
rect 9116 28430 9122 28436
rect 9478 28430 9484 28436
rect 9116 28390 9484 28430
rect 9116 28384 9122 28390
rect 9478 28384 9484 28390
rect 9536 28384 9542 28436
rect 4400 28290 4822 28350
rect 4880 28290 4886 28350
rect 4400 27900 4460 28290
rect 6420 28090 6480 28350
rect 8190 28340 8250 28346
rect 8190 28090 8250 28281
rect 23880 28220 23940 28226
rect 6420 28030 10242 28090
rect 10300 28030 10306 28090
rect 6420 27900 6480 28030
rect 4400 27840 6480 27900
rect 10100 27790 10160 28030
rect 11160 27890 11390 27950
rect 11450 27890 11456 27950
rect 11160 27790 11220 27890
rect 10100 27730 11220 27790
rect 16550 27100 16610 27106
rect 15490 26310 15550 26316
rect 15490 14778 15550 26250
rect 16550 15748 16610 27040
rect 23880 16718 23940 28160
rect 23880 16662 23882 16718
rect 23938 16662 23940 16718
rect 23880 16660 23940 16662
rect 23882 16653 23938 16660
rect 16550 15692 16552 15748
rect 16608 15692 16610 15748
rect 16550 15690 16610 15692
rect 16552 15683 16608 15690
rect 15490 14722 15492 14778
rect 15548 14722 15550 14778
rect 15490 14720 15550 14722
rect 15492 14713 15548 14720
<< via2 >>
rect 7012 35312 7068 35368
rect 6352 35222 6408 35278
rect 8502 34602 8558 34658
rect 8402 34422 8458 34478
rect 3792 34352 3848 34408
rect 3792 33982 3848 34038
rect 4212 33982 4268 34038
rect 7112 34112 7168 34168
rect 4012 33242 4068 33298
rect 10932 33102 10988 33158
rect 5952 32412 6008 32468
rect 7132 32372 7188 32428
rect 8982 31922 9038 31978
rect 7072 31302 7128 31358
rect 5582 31242 5638 31298
rect 7752 29422 7808 29478
rect 5942 29142 5998 29198
rect 11172 28812 11228 28868
rect 23882 16662 23938 16718
rect 16552 15692 16608 15748
rect 15492 14722 15548 14778
<< metal3 >>
rect 6330 35820 7550 35880
rect 6330 35550 6390 35820
rect 6050 35490 6770 35550
rect 6050 35280 6110 35490
rect 6710 35370 6770 35490
rect 7007 35370 7073 35373
rect 6710 35368 7073 35370
rect 6710 35312 7012 35368
rect 7068 35312 7073 35368
rect 6710 35310 7073 35312
rect 7007 35307 7073 35310
rect 6347 35280 6413 35283
rect 4210 35278 6413 35280
rect 4210 35222 6352 35278
rect 6408 35222 6413 35278
rect 4210 35220 6413 35222
rect 3787 34410 3853 34413
rect 2110 34408 3853 34410
rect 2110 34352 3792 34408
rect 3848 34352 3853 34408
rect 2110 34350 3853 34352
rect 194 33810 200 34210
rect 600 34040 606 34210
rect 1362 34040 1368 34042
rect 600 33980 1368 34040
rect 600 33810 606 33980
rect 1362 33978 1368 33980
rect 1432 33978 1438 34042
rect 2110 33630 2170 34350
rect 3787 34347 3853 34350
rect 2418 34042 2482 34048
rect 4210 34043 4270 35220
rect 6347 35217 6413 35220
rect 7490 35010 7550 35820
rect 7490 34950 8390 35010
rect 7490 34440 7550 34950
rect 8330 34900 8390 34950
rect 8330 34840 8920 34900
rect 8330 34660 8390 34840
rect 8497 34660 8563 34663
rect 8330 34658 8563 34660
rect 8330 34602 8502 34658
rect 8558 34602 8563 34658
rect 8330 34600 8563 34602
rect 8497 34597 8563 34600
rect 7240 34380 7550 34440
rect 8397 34480 8463 34483
rect 8860 34480 8920 34840
rect 8397 34478 8920 34480
rect 8397 34422 8402 34478
rect 8458 34422 8920 34478
rect 8397 34420 8920 34422
rect 8397 34417 8463 34420
rect 7107 34170 7173 34173
rect 7240 34170 7300 34380
rect 7107 34168 7300 34170
rect 7107 34112 7112 34168
rect 7168 34112 7300 34168
rect 7107 34110 7300 34112
rect 7107 34107 7173 34110
rect 3787 34040 3853 34043
rect 2482 34038 3853 34040
rect 2482 33982 3792 34038
rect 3848 33982 3853 34038
rect 2482 33980 3853 33982
rect 2418 33972 2482 33978
rect 3350 33700 3410 33980
rect 3787 33977 3853 33980
rect 4207 34038 4273 34043
rect 4207 33982 4212 34038
rect 4268 33982 4273 34038
rect 4207 33977 4273 33982
rect 3350 33640 4840 33700
rect 2110 33570 2810 33630
rect 794 33070 800 33470
rect 1200 33300 1206 33470
rect 2750 33300 2810 33570
rect 4007 33300 4073 33303
rect 1200 33298 4073 33300
rect 1200 33242 4012 33298
rect 4068 33242 4073 33298
rect 1200 33240 4073 33242
rect 1200 33070 1206 33240
rect 4007 33237 4073 33240
rect 4780 32470 4840 33640
rect 8550 33370 10990 33430
rect 8550 32640 8610 33370
rect 10930 33163 10990 33370
rect 10927 33158 10993 33163
rect 10927 33102 10932 33158
rect 10988 33102 10993 33158
rect 10927 33097 10993 33102
rect 5790 32580 9040 32640
rect 5790 32470 5850 32580
rect 5947 32470 6013 32473
rect 4780 32468 6013 32470
rect 4780 32412 5952 32468
rect 6008 32412 6013 32468
rect 7130 32433 7190 32580
rect 4780 32410 6013 32412
rect 5580 31480 5640 32410
rect 5947 32407 6013 32410
rect 7127 32428 7193 32433
rect 7127 32372 7132 32428
rect 7188 32372 7193 32428
rect 7127 32367 7193 32372
rect 8980 31983 9040 32580
rect 8977 31978 9043 31983
rect 8977 31922 8982 31978
rect 9038 31922 9043 31978
rect 8977 31917 9043 31922
rect 6180 31510 7130 31570
rect 6180 31480 6240 31510
rect 5310 31420 6240 31480
rect 5310 29830 5370 31420
rect 5580 31303 5640 31420
rect 7070 31363 7130 31510
rect 7067 31358 7133 31363
rect 5577 31298 5643 31303
rect 5577 31242 5582 31298
rect 5638 31242 5643 31298
rect 7067 31302 7072 31358
rect 7128 31302 7133 31358
rect 7067 31297 7133 31302
rect 5577 31237 5643 31242
rect 6390 30220 8890 30280
rect 6390 29830 6450 30220
rect 5310 29770 6760 29830
rect 5310 29440 5370 29770
rect 6700 29480 6760 29770
rect 7747 29480 7813 29483
rect 6700 29478 7813 29480
rect 5310 29380 6000 29440
rect 6700 29422 7752 29478
rect 7808 29422 7813 29478
rect 6700 29420 7813 29422
rect 7747 29417 7813 29420
rect 5940 29203 6000 29380
rect 8830 29350 8890 30220
rect 8830 29290 11230 29350
rect 5937 29198 6003 29203
rect 5937 29142 5942 29198
rect 5998 29142 6003 29198
rect 5937 29137 6003 29142
rect 11170 28873 11230 29290
rect 11167 28868 11233 28873
rect 11167 28812 11172 28868
rect 11228 28812 11233 28868
rect 11167 28807 11233 28812
rect 23877 16720 23943 16723
rect 23877 16718 29780 16720
rect 23877 16662 23882 16718
rect 23938 16662 29780 16718
rect 23877 16660 29780 16662
rect 23877 16657 23943 16660
rect 16547 15750 16613 15753
rect 16547 15748 25750 15750
rect 16547 15692 16552 15748
rect 16608 15692 25750 15748
rect 16547 15690 25750 15692
rect 16547 15687 16613 15690
rect 15487 14780 15553 14783
rect 15487 14778 21980 14780
rect 15487 14722 15492 14778
rect 15548 14722 21980 14778
rect 15487 14720 21980 14722
rect 15487 14717 15553 14720
rect 21920 720 21980 14720
rect 21920 660 22250 720
rect 22190 340 22250 660
rect 25690 390 25750 15690
rect 29720 800 29780 16660
rect 29720 740 30480 800
rect 22190 280 22750 340
rect 25690 330 26620 390
rect 22690 206 22750 280
rect 22630 200 22810 206
rect 26560 196 26620 330
rect 30420 196 30480 740
rect 22630 14 22810 20
rect 26500 190 26680 196
rect 26500 4 26680 10
rect 30360 190 30540 196
rect 30360 4 30540 10
<< via3 >>
rect 200 33810 600 34210
rect 1368 33978 1432 34042
rect 2418 33978 2482 34042
rect 800 33070 1200 33470
rect 22630 20 22810 200
rect 26500 10 26680 190
rect 30360 10 30540 190
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 34211 600 44152
rect 199 34210 601 34211
rect 199 33810 200 34210
rect 600 33810 601 34210
rect 199 33809 601 33810
rect 200 1000 600 33809
rect 800 33471 1200 44152
rect 1367 34042 1433 34043
rect 1367 33978 1368 34042
rect 1432 34040 1433 34042
rect 2417 34042 2483 34043
rect 2417 34040 2418 34042
rect 1432 33980 2418 34040
rect 1432 33978 1433 33980
rect 1367 33977 1433 33978
rect 2417 33978 2418 33980
rect 2482 33978 2483 34042
rect 2417 33977 2483 33978
rect 799 33470 1201 33471
rect 799 33070 800 33470
rect 1200 33070 1201 33470
rect 799 33069 1201 33070
rect 800 1000 1200 33069
rect 22629 200 22811 201
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22629 20 22630 200
rect 22810 20 22814 200
rect 22629 19 22814 20
rect 22634 0 22814 19
rect 26498 191 26678 200
rect 30362 191 30542 200
rect 26498 190 26681 191
rect 26498 10 26500 190
rect 26680 10 26681 190
rect 26498 9 26681 10
rect 30359 190 30542 191
rect 30359 10 30360 190
rect 30540 10 30542 190
rect 30359 9 30542 10
rect 26498 0 26678 9
rect 30362 0 30542 9
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4670 0 1 28450
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_1
timestamp 1723858470
transform 1 0 10380 0 1 28080
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6340 0 1 34510
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1723858470
transform 1 0 6250 0 1 33450
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1723858470
transform 1 0 6040 0 1 31680
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1723858470
transform 1 0 6048 0 1 30708
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1723858470
transform 1 0 7528 0 1 28498
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7860 0 1 33910
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1723858470
transform 1 0 8010 0 1 31180
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7128 0 1 34508
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1723858470
transform 1 0 6908 0 1 33448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1723858470
transform 1 0 6738 0 1 31688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1723858470
transform 1 0 6708 0 1 30708
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1723858470
transform 1 0 8650 0 1 33850
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1723858470
transform 1 0 8788 0 1 31178
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1723858470
transform 1 0 11308 0 1 32178
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1723858470
transform 1 0 8178 0 1 28488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1723858470
transform 1 0 5708 0 1 28458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1723858470
transform 1 0 11378 0 1 28078
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10138 0 1 32188
box -38 -48 682 592
<< labels >>
rlabel metal4 s 28766 44952 28826 45152 6 clk
port 0 nsew default input
rlabel metal4 s 29318 44952 29378 45152 6 ena
port 1 nsew default input
rlabel metal4 s 28214 44952 28274 45152 6 rst_n
port 2 nsew default input
rlabel metal4 s 30362 0 30542 200 6 ua[0]
port 3 nsew default bidirectional
rlabel metal4 s 26498 0 26678 200 6 ua[1]
port 4 nsew default bidirectional
rlabel metal4 s 22634 0 22814 200 6 ua[2]
port 5 nsew default bidirectional
rlabel metal4 s 18770 0 18950 200 6 ua[3]
port 6 nsew default bidirectional
rlabel metal4 s 14906 0 15086 200 6 ua[4]
port 7 nsew default bidirectional
rlabel metal4 s 11042 0 11222 200 6 ua[5]
port 8 nsew default bidirectional
rlabel metal4 s 7178 0 7358 200 6 ua[6]
port 9 nsew default bidirectional
rlabel metal4 s 3314 0 3494 200 6 ua[7]
port 10 nsew default bidirectional
rlabel metal4 s 27662 44952 27722 45152 6 ui_in[0]
port 11 nsew default input
rlabel metal4 s 27110 44952 27170 45152 6 ui_in[1]
port 12 nsew default input
rlabel metal4 s 26558 44952 26618 45152 6 ui_in[2]
port 13 nsew default input
rlabel metal4 s 26006 44952 26066 45152 6 ui_in[3]
port 14 nsew default input
rlabel metal4 s 25454 44952 25514 45152 6 ui_in[4]
port 15 nsew default input
rlabel metal4 s 24902 44952 24962 45152 6 ui_in[5]
port 16 nsew default input
rlabel metal4 s 24350 44952 24410 45152 6 ui_in[6]
port 17 nsew default input
rlabel metal4 s 23798 44952 23858 45152 6 ui_in[7]
port 18 nsew default input
rlabel metal4 s 23246 44952 23306 45152 6 uio_in[0]
port 19 nsew default input
rlabel metal4 s 22694 44952 22754 45152 6 uio_in[1]
port 20 nsew default input
rlabel metal4 s 22142 44952 22202 45152 6 uio_in[2]
port 21 nsew default input
rlabel metal4 s 21590 44952 21650 45152 6 uio_in[3]
port 22 nsew default input
rlabel metal4 s 21038 44952 21098 45152 6 uio_in[4]
port 23 nsew default input
rlabel metal4 s 20486 44952 20546 45152 6 uio_in[5]
port 24 nsew default input
rlabel metal4 s 19934 44952 19994 45152 6 uio_in[6]
port 25 nsew default input
rlabel metal4 s 19382 44952 19442 45152 6 uio_in[7]
port 26 nsew default input
rlabel metal4 s 9998 44952 10058 45152 6 uio_oe[0]
port 27 nsew default tristate
rlabel metal4 s 9446 44952 9506 45152 6 uio_oe[1]
port 28 nsew default tristate
rlabel metal4 s 8894 44952 8954 45152 6 uio_oe[2]
port 29 nsew default tristate
rlabel metal4 s 8342 44952 8402 45152 6 uio_oe[3]
port 30 nsew default tristate
rlabel metal4 s 7790 44952 7850 45152 6 uio_oe[4]
port 31 nsew default tristate
rlabel metal4 s 7238 44952 7298 45152 6 uio_oe[5]
port 32 nsew default tristate
rlabel metal4 s 6686 44952 6746 45152 6 uio_oe[6]
port 33 nsew default tristate
rlabel metal4 s 6134 44952 6194 45152 6 uio_oe[7]
port 34 nsew default tristate
rlabel metal4 s 14414 44952 14474 45152 6 uio_out[0]
port 35 nsew default tristate
rlabel metal4 s 13862 44952 13922 45152 6 uio_out[1]
port 36 nsew default tristate
rlabel metal4 s 13310 44952 13370 45152 6 uio_out[2]
port 37 nsew default tristate
rlabel metal4 s 12758 44952 12818 45152 6 uio_out[3]
port 38 nsew default tristate
rlabel metal4 s 12206 44952 12266 45152 6 uio_out[4]
port 39 nsew default tristate
rlabel metal4 s 11654 44952 11714 45152 6 uio_out[5]
port 40 nsew default tristate
rlabel metal4 s 11102 44952 11162 45152 6 uio_out[6]
port 41 nsew default tristate
rlabel metal4 s 10550 44952 10610 45152 6 uio_out[7]
port 42 nsew default tristate
rlabel metal4 s 18830 44952 18890 45152 6 uo_out[0]
port 43 nsew default tristate
rlabel metal4 s 18278 44952 18338 45152 6 uo_out[1]
port 44 nsew default tristate
rlabel metal4 s 17726 44952 17786 45152 6 uo_out[2]
port 45 nsew default tristate
rlabel metal4 s 17174 44952 17234 45152 6 uo_out[3]
port 46 nsew default tristate
rlabel metal4 s 16622 44952 16682 45152 6 uo_out[4]
port 47 nsew default tristate
rlabel metal4 s 16070 44952 16130 45152 6 uo_out[5]
port 48 nsew default tristate
rlabel metal4 s 15518 44952 15578 45152 6 uo_out[6]
port 49 nsew default tristate
rlabel metal4 s 14966 44952 15026 45152 6 uo_out[7]
port 50 nsew default tristate
flabel metal4 200 1000 600 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< end >>
