VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_17
  CLASS BLOCK ;
  FOREIGN tt_um_test_17 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 142.860 224.760 143.160 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 145.620 224.760 145.920 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 140.100 224.760 140.400 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 52.550 142.525 53.145 142.865 ;
        RECT 52.550 141.205 52.725 142.525 ;
        RECT 52.550 141.100 53.145 141.205 ;
        RECT 52.550 140.800 53.930 141.100 ;
        RECT 52.550 140.655 53.145 140.800 ;
      LAYER met1 ;
        RECT 53.600 140.800 118.760 141.100 ;
      LAYER met2 ;
        RECT 118.430 83.300 118.730 141.130 ;
        RECT 118.440 83.265 118.720 83.300 ;
      LAYER met3 ;
        RECT 118.415 83.600 118.745 83.615 ;
        RECT 118.415 83.300 147.930 83.600 ;
        RECT 118.415 83.285 118.745 83.300 ;
        RECT 147.630 4.000 147.930 83.300 ;
        RECT 147.630 3.700 151.430 4.000 ;
        RECT 151.130 0.980 151.430 3.700 ;
        RECT 150.830 0.020 151.730 0.980 ;
      LAYER met4 ;
        RECT 150.840 0.955 151.740 1.000 ;
        RECT 150.825 0.045 151.740 0.955 ;
        RECT 150.840 0.000 151.740 0.045 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 29.550 159.700 29.880 159.715 ;
        RECT 28.380 159.500 29.880 159.700 ;
        RECT 29.550 159.475 29.880 159.500 ;
      LAYER met1 ;
        RECT 23.500 159.700 23.760 159.760 ;
        RECT 16.980 159.500 23.760 159.700 ;
        RECT 16.980 135.500 17.280 159.500 ;
        RECT 23.500 159.440 23.760 159.500 ;
        RECT 25.600 159.700 25.860 159.760 ;
        RECT 28.335 159.700 28.625 159.715 ;
        RECT 25.600 159.500 28.625 159.700 ;
        RECT 25.600 159.440 25.860 159.500 ;
        RECT 28.335 159.485 28.625 159.500 ;
        RECT 16.980 135.200 82.110 135.500 ;
      LAYER met2 ;
        RECT 23.470 159.700 23.790 159.730 ;
        RECT 25.570 159.700 25.890 159.730 ;
        RECT 23.470 159.500 25.890 159.700 ;
        RECT 23.470 159.470 23.790 159.500 ;
        RECT 25.570 159.470 25.890 159.500 ;
        RECT 81.780 78.450 82.080 135.530 ;
        RECT 81.790 78.415 82.070 78.450 ;
      LAYER met3 ;
        RECT 81.765 78.750 82.095 78.765 ;
        RECT 81.765 78.450 127.780 78.750 ;
        RECT 81.765 78.435 82.095 78.450 ;
        RECT 127.480 1.950 127.780 78.450 ;
        RECT 127.480 1.650 132.130 1.950 ;
        RECT 131.830 0.980 132.130 1.650 ;
        RECT 131.530 0.020 132.430 0.980 ;
      LAYER met4 ;
        RECT 131.520 0.955 132.420 1.000 ;
        RECT 131.520 0.045 132.435 0.955 ;
        RECT 131.520 0.000 132.420 0.045 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 31.050 173.850 31.380 173.865 ;
        RECT 30.030 173.650 31.380 173.850 ;
        RECT 31.050 173.625 31.380 173.650 ;
      LAYER met1 ;
        RECT 29.985 173.850 30.275 173.865 ;
        RECT 13.780 173.650 30.275 173.850 ;
        RECT 13.780 131.550 14.080 173.650 ;
        RECT 29.985 173.635 30.275 173.650 ;
        RECT 13.780 131.250 76.810 131.550 ;
      LAYER met2 ;
        RECT 76.480 73.600 76.780 131.580 ;
        RECT 76.490 73.565 76.770 73.600 ;
      LAYER met3 ;
        RECT 76.465 73.900 76.795 73.915 ;
        RECT 76.465 73.600 108.930 73.900 ;
        RECT 76.465 73.585 76.795 73.600 ;
        RECT 108.630 3.600 108.930 73.600 ;
        RECT 108.630 3.300 110.280 3.600 ;
        RECT 109.980 1.700 110.280 3.300 ;
        RECT 109.980 1.400 112.780 1.700 ;
        RECT 112.480 1.030 112.780 1.400 ;
        RECT 112.180 0.070 113.080 1.030 ;
      LAYER met4 ;
        RECT 112.175 1.000 113.085 1.005 ;
        RECT 112.175 0.095 113.100 1.000 ;
        RECT 112.200 0.000 113.100 0.095 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 92.880 0.000 93.780 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 73.560 0.000 74.460 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 54.240 0.000 55.140 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 34.920 0.000 35.820 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 15.600 0.000 16.500 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 137.340 224.760 137.640 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 134.580 224.760 134.880 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 131.820 224.760 132.120 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 129.060 224.760 129.360 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 126.300 224.760 126.600 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 123.540 224.760 123.840 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 120.780 224.760 121.080 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 118.020 224.760 118.320 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 115.260 224.760 115.560 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 112.500 224.760 112.800 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 109.740 224.760 110.040 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 106.980 224.760 107.280 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 104.220 224.760 104.520 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 101.460 224.760 101.760 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 98.700 224.760 99.000 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 95.940 224.760 96.240 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 49.020 224.760 49.320 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 46.260 224.760 46.560 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 43.500 224.760 43.800 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 40.740 224.760 41.040 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 37.980 224.760 38.280 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 35.220 224.760 35.520 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 32.460 224.760 32.760 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 29.700 224.760 30.000 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 71.100 224.760 71.400 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 68.340 224.760 68.640 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 65.580 224.760 65.880 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 62.820 224.760 63.120 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 60.060 224.760 60.360 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 57.300 224.760 57.600 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 54.540 224.760 54.840 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 51.780 224.760 52.080 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 93.180 224.760 93.480 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 90.420 224.760 90.720 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 87.660 224.760 87.960 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 84.900 224.760 85.200 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 82.140 224.760 82.440 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 79.380 224.760 79.680 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 76.620 224.760 76.920 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 73.860 224.760 74.160 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 30.540 175.450 33.580 175.460 ;
        RECT 30.540 173.855 35.320 175.450 ;
        RECT 33.560 173.845 35.320 173.855 ;
        RECT 38.140 172.160 41.180 172.460 ;
        RECT 38.140 170.855 42.930 172.160 ;
        RECT 41.160 170.555 42.930 170.855 ;
        RECT 30.090 170.150 32.680 170.160 ;
        RECT 30.090 168.555 34.220 170.150 ;
        RECT 32.660 168.545 34.220 168.555 ;
        RECT 49.530 163.800 54.430 163.850 ;
        RECT 49.530 162.245 56.220 163.800 ;
        RECT 54.360 162.195 56.220 162.245 ;
        RECT 31.660 161.310 33.370 161.350 ;
        RECT 29.040 159.745 33.370 161.310 ;
        RECT 29.040 159.705 31.780 159.745 ;
        RECT 38.890 158.800 41.930 158.810 ;
        RECT 38.890 157.205 43.620 158.800 ;
        RECT 41.910 157.195 43.620 157.205 ;
        RECT 29.080 154.845 33.220 156.450 ;
        RECT 36.480 145.350 39.080 145.400 ;
        RECT 26.560 145.160 28.220 145.200 ;
        RECT 22.190 143.595 28.220 145.160 ;
        RECT 36.480 143.795 40.570 145.350 ;
        RECT 38.910 143.745 40.570 143.795 ;
        RECT 22.190 143.555 26.580 143.595 ;
        RECT 50.740 143.300 54.830 143.310 ;
        RECT 50.740 141.705 56.570 143.300 ;
        RECT 54.810 141.695 56.570 141.705 ;
      LAYER li1 ;
        RECT 30.730 175.185 32.110 175.355 ;
        RECT 31.070 174.045 31.280 175.185 ;
        RECT 34.670 175.175 35.130 175.345 ;
        RECT 34.755 174.010 35.045 175.175 ;
        RECT 38.330 172.185 39.710 172.355 ;
        RECT 39.285 171.045 39.615 172.185 ;
        RECT 42.280 171.885 42.740 172.055 ;
        RECT 42.365 170.720 42.655 171.885 ;
        RECT 30.280 169.885 31.660 170.055 ;
        RECT 30.620 168.745 30.830 169.885 ;
        RECT 33.570 169.875 34.030 170.045 ;
        RECT 33.655 168.710 33.945 169.875 ;
        RECT 49.720 163.575 52.940 163.745 ;
        RECT 50.775 162.725 50.945 163.575 ;
        RECT 51.615 163.065 51.785 163.575 ;
        RECT 55.570 163.525 56.030 163.695 ;
        RECT 55.655 162.360 55.945 163.525 ;
        RECT 29.230 161.035 30.610 161.205 ;
        RECT 32.720 161.075 33.180 161.245 ;
        RECT 29.570 159.895 29.780 161.035 ;
        RECT 32.805 159.910 33.095 161.075 ;
        RECT 39.080 158.535 40.460 158.705 ;
        RECT 40.035 157.395 40.365 158.535 ;
        RECT 42.970 158.525 43.430 158.695 ;
        RECT 43.055 157.360 43.345 158.525 ;
        RECT 29.270 156.175 30.650 156.345 ;
        RECT 32.570 156.175 33.030 156.345 ;
        RECT 29.610 155.035 29.820 156.175 ;
        RECT 32.655 155.010 32.945 156.175 ;
        RECT 36.670 145.125 38.050 145.295 ;
        RECT 22.380 144.885 24.680 145.055 ;
        RECT 27.570 144.925 28.030 145.095 ;
        RECT 22.895 144.485 23.830 144.885 ;
        RECT 27.655 143.760 27.945 144.925 ;
        RECT 37.010 143.985 37.220 145.125 ;
        RECT 39.920 145.075 40.380 145.245 ;
        RECT 40.005 143.910 40.295 145.075 ;
        RECT 50.930 143.035 53.230 143.205 ;
        RECT 51.445 142.635 52.380 143.035 ;
        RECT 55.920 143.025 56.380 143.195 ;
        RECT 56.005 141.860 56.295 143.025 ;
      LAYER met1 ;
        RECT 31.490 176.395 31.780 176.430 ;
        RECT 31.490 176.070 31.795 176.395 ;
        RECT 31.505 175.510 31.795 176.070 ;
        RECT 30.730 175.030 32.110 175.510 ;
        RECT 34.730 175.500 35.030 176.880 ;
        RECT 34.670 175.020 35.130 175.500 ;
        RECT 42.380 173.300 42.680 173.330 ;
        RECT 42.375 172.970 42.680 173.300 ;
        RECT 38.330 172.400 39.710 172.510 ;
        RECT 40.130 172.400 40.430 172.430 ;
        RECT 38.330 172.100 40.430 172.400 ;
        RECT 42.375 172.210 42.675 172.970 ;
        RECT 38.330 172.030 39.710 172.100 ;
        RECT 40.130 172.070 40.430 172.100 ;
        RECT 42.280 171.730 42.740 172.210 ;
        RECT 28.235 170.655 30.885 170.945 ;
        RECT 23.940 170.195 24.230 170.230 ;
        RECT 28.235 170.195 28.525 170.655 ;
        RECT 30.595 170.210 30.885 170.655 ;
        RECT 23.935 169.905 28.525 170.195 ;
        RECT 23.940 169.870 24.230 169.905 ;
        RECT 30.280 169.730 31.660 170.210 ;
        RECT 33.630 170.200 33.925 170.880 ;
        RECT 33.570 169.720 34.030 170.200 ;
        RECT 54.780 164.895 55.930 164.900 ;
        RECT 51.415 164.605 55.930 164.895 ;
        RECT 51.415 163.900 51.705 164.605 ;
        RECT 53.650 164.600 54.010 164.605 ;
        RECT 54.780 164.595 55.930 164.605 ;
        RECT 49.720 163.420 52.940 163.900 ;
        RECT 55.625 163.850 55.930 164.595 ;
        RECT 55.570 163.370 56.030 163.850 ;
        RECT 29.540 162.345 29.830 162.380 ;
        RECT 29.540 162.020 29.835 162.345 ;
        RECT 33.630 162.145 33.925 162.180 ;
        RECT 29.545 161.360 29.835 162.020 ;
        RECT 32.780 161.850 33.925 162.145 ;
        RECT 32.780 161.400 33.075 161.850 ;
        RECT 33.630 161.820 33.925 161.850 ;
        RECT 29.230 160.880 30.610 161.360 ;
        RECT 32.720 160.920 33.180 161.400 ;
        RECT 43.030 159.900 43.330 159.930 ;
        RECT 39.530 159.895 43.330 159.900 ;
        RECT 39.395 159.600 43.330 159.895 ;
        RECT 39.395 158.860 39.685 159.600 ;
        RECT 39.080 158.380 40.460 158.860 ;
        RECT 43.030 158.850 43.330 159.600 ;
        RECT 42.970 158.370 43.430 158.850 ;
        RECT 33.530 156.800 33.830 156.830 ;
        RECT 28.090 156.500 28.380 156.530 ;
        RECT 32.680 156.500 33.830 156.800 ;
        RECT 28.085 156.210 30.650 156.500 ;
        RECT 28.090 156.170 28.380 156.210 ;
        RECT 29.270 156.020 30.650 156.210 ;
        RECT 32.570 156.020 33.030 156.500 ;
        RECT 33.530 156.470 33.830 156.500 ;
        RECT 37.750 146.400 38.115 146.405 ;
        RECT 37.030 146.395 40.280 146.400 ;
        RECT 36.985 146.095 40.280 146.395 ;
        RECT 27.680 146.000 27.985 146.035 ;
        RECT 27.675 145.995 27.985 146.000 ;
        RECT 23.155 145.705 27.985 145.995 ;
        RECT 23.155 145.210 23.445 145.705 ;
        RECT 27.675 145.670 27.985 145.705 ;
        RECT 27.675 145.250 27.980 145.670 ;
        RECT 36.985 145.450 37.275 146.095 ;
        RECT 22.380 144.730 24.680 145.210 ;
        RECT 27.570 144.770 28.030 145.250 ;
        RECT 36.670 144.970 38.050 145.450 ;
        RECT 39.975 145.400 40.280 146.095 ;
        RECT 39.920 144.920 40.380 145.400 ;
        RECT 52.180 144.345 52.470 144.380 ;
        RECT 52.165 144.020 52.470 144.345 ;
        RECT 52.165 143.360 52.455 144.020 ;
        RECT 50.930 142.880 53.230 143.360 ;
        RECT 55.980 143.350 56.280 144.380 ;
        RECT 55.920 142.870 56.380 143.350 ;
      LAYER met2 ;
        RECT 34.090 176.850 34.370 176.885 ;
        RECT 34.080 176.550 35.060 176.850 ;
        RECT 34.090 176.515 34.370 176.550 ;
        RECT 30.790 176.400 31.070 176.435 ;
        RECT 30.780 176.100 31.810 176.400 ;
        RECT 30.790 176.065 31.070 176.100 ;
        RECT 41.540 173.300 41.820 173.335 ;
        RECT 41.530 173.000 42.710 173.300 ;
        RECT 41.540 172.965 41.820 173.000 ;
        RECT 41.040 172.400 41.320 172.435 ;
        RECT 40.100 172.100 41.320 172.400 ;
        RECT 41.040 172.065 41.320 172.100 ;
        RECT 34.590 170.850 34.870 170.885 ;
        RECT 33.600 170.550 34.880 170.850 ;
        RECT 34.590 170.515 34.870 170.550 ;
        RECT 17.990 170.200 18.270 170.235 ;
        RECT 17.980 169.900 24.260 170.200 ;
        RECT 17.990 169.865 18.270 169.900 ;
        RECT 53.680 165.790 53.980 165.800 ;
        RECT 53.645 165.510 54.015 165.790 ;
        RECT 53.680 164.570 53.980 165.510 ;
        RECT 28.790 162.350 29.070 162.385 ;
        RECT 28.780 162.050 29.860 162.350 ;
        RECT 33.600 162.140 34.980 162.150 ;
        RECT 28.790 162.015 29.070 162.050 ;
        RECT 33.600 161.860 35.015 162.140 ;
        RECT 33.600 161.850 34.980 161.860 ;
        RECT 43.000 159.890 44.230 159.900 ;
        RECT 43.000 159.610 44.265 159.890 ;
        RECT 43.000 159.600 44.230 159.610 ;
        RECT 33.500 156.790 34.680 156.800 ;
        RECT 33.500 156.510 34.715 156.790 ;
        RECT 33.500 156.500 34.680 156.510 ;
        RECT 26.930 156.490 28.410 156.500 ;
        RECT 26.895 156.210 28.410 156.490 ;
        RECT 26.930 156.200 28.410 156.210 ;
        RECT 37.790 147.400 38.070 147.435 ;
        RECT 37.780 146.435 38.080 147.400 ;
        RECT 37.780 146.070 38.085 146.435 ;
        RECT 27.650 146.000 28.015 146.005 ;
        RECT 27.650 145.990 29.030 146.000 ;
        RECT 27.650 145.710 29.065 145.990 ;
        RECT 27.650 145.700 29.030 145.710 ;
        RECT 52.150 144.050 56.310 144.350 ;
      LAYER met3 ;
        RECT 30.680 179.100 36.780 179.400 ;
        RECT 30.680 177.750 30.980 179.100 ;
        RECT 29.280 177.450 32.880 177.750 ;
        RECT 29.280 176.400 29.580 177.450 ;
        RECT 32.580 176.850 32.880 177.450 ;
        RECT 34.065 176.850 34.395 176.865 ;
        RECT 32.580 176.550 34.395 176.850 ;
        RECT 34.065 176.535 34.395 176.550 ;
        RECT 30.765 176.400 31.095 176.415 ;
        RECT 20.080 176.100 31.095 176.400 ;
        RECT 0.000 170.200 2.060 171.050 ;
        RECT 5.840 170.200 6.220 170.210 ;
        RECT 0.000 169.900 6.220 170.200 ;
        RECT 0.000 169.050 2.060 169.900 ;
        RECT 5.840 169.890 6.220 169.900 ;
        RECT 11.120 170.200 11.440 170.240 ;
        RECT 20.080 170.215 20.380 176.100 ;
        RECT 30.765 176.085 31.095 176.100 ;
        RECT 36.480 175.050 36.780 179.100 ;
        RECT 36.480 174.750 40.980 175.050 ;
        RECT 36.480 172.200 36.780 174.750 ;
        RECT 40.680 174.500 40.980 174.750 ;
        RECT 40.680 174.200 43.630 174.500 ;
        RECT 40.680 173.300 40.980 174.200 ;
        RECT 41.515 173.300 41.845 173.315 ;
        RECT 40.680 173.000 41.845 173.300 ;
        RECT 41.515 172.985 41.845 173.000 ;
        RECT 35.230 171.900 36.780 172.200 ;
        RECT 41.015 172.400 41.345 172.415 ;
        RECT 43.330 172.400 43.630 174.200 ;
        RECT 41.015 172.100 43.630 172.400 ;
        RECT 41.015 172.085 41.345 172.100 ;
        RECT 34.565 170.850 34.895 170.865 ;
        RECT 35.230 170.850 35.530 171.900 ;
        RECT 34.565 170.550 35.530 170.850 ;
        RECT 34.565 170.535 34.895 170.550 ;
        RECT 17.965 170.200 18.295 170.215 ;
        RECT 11.120 169.900 18.295 170.200 ;
        RECT 11.120 169.860 11.440 169.900 ;
        RECT 15.780 168.500 16.080 169.900 ;
        RECT 17.965 169.885 18.295 169.900 ;
        RECT 20.065 169.885 20.395 170.215 ;
        RECT 15.780 168.200 23.230 168.500 ;
        RECT 22.930 162.350 23.230 168.200 ;
        RECT 41.780 166.850 53.980 167.150 ;
        RECT 41.780 163.200 42.080 166.850 ;
        RECT 53.680 165.815 53.980 166.850 ;
        RECT 53.665 165.485 53.995 165.815 ;
        RECT 27.980 162.900 44.230 163.200 ;
        RECT 27.980 162.350 28.280 162.900 ;
        RECT 28.765 162.350 29.095 162.365 ;
        RECT 22.930 162.050 29.095 162.350 ;
        RECT 34.680 162.165 34.980 162.900 ;
        RECT 26.930 157.400 27.230 162.050 ;
        RECT 28.765 162.035 29.095 162.050 ;
        RECT 34.665 161.835 34.995 162.165 ;
        RECT 43.930 159.915 44.230 162.900 ;
        RECT 43.915 159.585 44.245 159.915 ;
        RECT 29.930 157.550 34.680 157.850 ;
        RECT 29.930 157.400 30.230 157.550 ;
        RECT 25.580 157.100 30.230 157.400 ;
        RECT 25.580 149.150 25.880 157.100 ;
        RECT 26.930 156.515 27.230 157.100 ;
        RECT 34.380 156.815 34.680 157.550 ;
        RECT 26.915 156.185 27.245 156.515 ;
        RECT 34.365 156.485 34.695 156.815 ;
        RECT 30.980 151.100 43.480 151.400 ;
        RECT 30.980 149.150 31.280 151.100 ;
        RECT 25.580 148.850 32.830 149.150 ;
        RECT 25.580 147.200 25.880 148.850 ;
        RECT 32.530 147.400 32.830 148.850 ;
        RECT 37.765 147.400 38.095 147.415 ;
        RECT 25.580 146.900 29.030 147.200 ;
        RECT 32.530 147.100 38.095 147.400 ;
        RECT 37.765 147.085 38.095 147.100 ;
        RECT 28.730 146.015 29.030 146.900 ;
        RECT 43.180 146.750 43.480 151.100 ;
        RECT 43.180 146.450 55.180 146.750 ;
        RECT 28.715 145.685 29.045 146.015 ;
        RECT 54.880 144.365 55.180 146.450 ;
        RECT 54.865 144.035 55.195 144.365 ;
      LAYER met4 ;
        RECT 0.030 171.055 2.030 220.760 ;
        RECT 0.025 169.045 2.035 171.055 ;
        RECT 5.865 170.200 6.195 170.215 ;
        RECT 11.115 170.200 11.445 170.215 ;
        RECT 5.865 169.900 11.445 170.200 ;
        RECT 5.865 169.885 6.195 169.900 ;
        RECT 11.115 169.885 11.445 169.900 ;
        RECT 0.030 5.000 2.030 169.045 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 34.685 172.730 35.115 173.515 ;
        RECT 42.295 169.440 42.725 170.225 ;
        RECT 33.585 167.430 34.015 168.215 ;
        RECT 55.585 161.080 56.015 161.865 ;
        RECT 32.735 158.630 33.165 159.415 ;
        RECT 42.985 156.080 43.415 156.865 ;
        RECT 32.585 153.730 33.015 154.515 ;
        RECT 27.585 142.480 28.015 143.265 ;
        RECT 39.935 142.630 40.365 143.415 ;
        RECT 55.935 140.580 56.365 141.365 ;
      LAYER li1 ;
        RECT 31.050 172.635 31.280 173.455 ;
        RECT 30.730 172.465 32.110 172.635 ;
        RECT 34.755 172.625 35.045 173.350 ;
        RECT 34.670 172.455 35.130 172.625 ;
        RECT 38.435 169.635 38.675 170.445 ;
        RECT 39.345 169.635 39.615 170.445 ;
        RECT 38.330 169.465 39.710 169.635 ;
        RECT 42.365 169.335 42.655 170.060 ;
        RECT 42.280 169.165 42.740 169.335 ;
        RECT 30.600 167.335 30.830 168.155 ;
        RECT 30.280 167.165 31.660 167.335 ;
        RECT 33.655 167.325 33.945 168.050 ;
        RECT 33.570 167.155 34.030 167.325 ;
        RECT 49.855 161.025 50.185 161.415 ;
        RECT 50.695 161.025 51.025 161.415 ;
        RECT 52.565 161.025 52.855 161.860 ;
        RECT 49.720 160.855 52.940 161.025 ;
        RECT 55.655 160.975 55.945 161.700 ;
        RECT 55.570 160.805 56.030 160.975 ;
        RECT 29.550 158.485 29.780 159.305 ;
        RECT 32.805 158.525 33.095 159.250 ;
        RECT 29.230 158.315 30.610 158.485 ;
        RECT 32.720 158.355 33.180 158.525 ;
        RECT 39.185 155.985 39.425 156.795 ;
        RECT 40.095 155.985 40.365 156.795 ;
        RECT 39.080 155.815 40.460 155.985 ;
        RECT 43.055 155.975 43.345 156.700 ;
        RECT 42.970 155.805 43.430 155.975 ;
        RECT 29.590 153.625 29.820 154.445 ;
        RECT 32.655 153.625 32.945 154.350 ;
        RECT 29.270 153.455 30.650 153.625 ;
        RECT 32.570 153.455 33.030 153.625 ;
        RECT 22.895 142.335 23.830 142.735 ;
        RECT 27.655 142.375 27.945 143.100 ;
        RECT 36.990 142.575 37.220 143.395 ;
        RECT 36.670 142.405 38.050 142.575 ;
        RECT 40.005 142.525 40.295 143.250 ;
        RECT 22.380 142.165 24.680 142.335 ;
        RECT 27.570 142.205 28.030 142.375 ;
        RECT 39.920 142.355 40.380 142.525 ;
        RECT 51.445 140.485 52.380 140.885 ;
        RECT 50.930 140.315 53.230 140.485 ;
        RECT 56.005 140.475 56.295 141.200 ;
        RECT 55.920 140.305 56.380 140.475 ;
      LAYER met1 ;
        RECT 30.730 172.310 32.110 172.790 ;
        RECT 23.890 172.045 24.180 172.080 ;
        RECT 31.045 172.045 31.335 172.310 ;
        RECT 34.670 172.300 35.130 172.780 ;
        RECT 23.885 171.755 31.335 172.045 ;
        RECT 34.780 171.770 35.080 172.300 ;
        RECT 23.890 171.720 24.180 171.755 ;
        RECT 37.690 169.600 37.980 169.630 ;
        RECT 38.330 169.600 39.710 169.790 ;
        RECT 37.685 169.310 39.710 169.600 ;
        RECT 37.690 169.270 37.980 169.310 ;
        RECT 42.280 169.010 42.740 169.490 ;
        RECT 42.330 168.270 42.630 169.010 ;
        RECT 30.280 167.010 31.660 167.490 ;
        RECT 25.690 166.495 25.980 166.530 ;
        RECT 30.595 166.495 30.885 167.010 ;
        RECT 33.570 167.000 34.030 167.480 ;
        RECT 25.685 166.205 30.885 166.495 ;
        RECT 33.625 166.680 33.925 167.000 ;
        RECT 33.625 166.350 33.930 166.680 ;
        RECT 33.630 166.320 33.930 166.350 ;
        RECT 25.690 166.170 25.980 166.205 ;
        RECT 48.790 160.990 49.080 161.030 ;
        RECT 49.720 160.990 52.940 161.180 ;
        RECT 48.785 160.700 52.940 160.990 ;
        RECT 48.790 160.670 49.080 160.700 ;
        RECT 55.570 160.650 56.030 161.130 ;
        RECT 55.630 159.720 55.930 160.650 ;
        RECT 29.230 158.160 30.610 158.640 ;
        RECT 32.720 158.250 33.180 158.680 ;
        RECT 33.630 158.250 33.930 158.280 ;
        RECT 32.720 158.200 33.930 158.250 ;
        RECT 25.590 157.845 25.880 157.880 ;
        RECT 29.545 157.845 29.835 158.160 ;
        RECT 32.775 157.950 33.930 158.200 ;
        RECT 33.630 157.920 33.930 157.950 ;
        RECT 25.585 157.555 29.835 157.845 ;
        RECT 25.590 157.520 25.880 157.555 ;
        RECT 38.290 155.950 38.580 155.980 ;
        RECT 39.080 155.950 40.460 156.140 ;
        RECT 38.285 155.660 40.460 155.950 ;
        RECT 38.290 155.620 38.580 155.660 ;
        RECT 42.970 155.650 43.430 156.130 ;
        RECT 43.075 155.085 43.380 155.650 ;
        RECT 43.075 154.750 43.385 155.085 ;
        RECT 43.080 154.720 43.385 154.750 ;
        RECT 29.270 153.300 30.650 153.780 ;
        RECT 32.570 153.300 33.030 153.780 ;
        RECT 29.585 153.130 29.875 153.300 ;
        RECT 29.585 152.805 29.880 153.130 ;
        RECT 29.590 152.770 29.880 152.805 ;
        RECT 32.630 152.600 32.930 153.300 ;
        RECT 32.600 152.300 32.960 152.600 ;
        RECT 35.890 142.540 36.180 142.580 ;
        RECT 36.670 142.540 38.050 142.730 ;
        RECT 22.380 142.010 24.680 142.490 ;
        RECT 27.570 142.050 28.030 142.530 ;
        RECT 35.885 142.250 38.050 142.540 ;
        RECT 35.890 142.220 36.180 142.250 ;
        RECT 39.920 142.200 40.380 142.680 ;
        RECT 28.480 142.050 28.780 142.080 ;
        RECT 23.155 141.780 23.445 142.010 ;
        RECT 23.140 141.455 23.445 141.780 ;
        RECT 27.630 141.750 28.780 142.050 ;
        RECT 39.980 141.950 40.280 142.200 ;
        RECT 28.480 141.720 28.780 141.750 ;
        RECT 39.985 141.700 40.280 141.950 ;
        RECT 23.140 141.420 23.430 141.455 ;
        RECT 39.950 141.405 40.310 141.700 ;
        RECT 50.240 140.450 50.530 140.480 ;
        RECT 50.930 140.450 53.230 140.640 ;
        RECT 50.235 140.160 53.230 140.450 ;
        RECT 50.240 140.120 50.530 140.160 ;
        RECT 55.920 140.150 56.380 140.630 ;
        RECT 55.980 139.420 56.280 140.150 ;
      LAYER met2 ;
        RECT 17.990 172.050 18.270 172.085 ;
        RECT 17.980 171.750 24.210 172.050 ;
        RECT 31.580 171.800 35.110 172.100 ;
        RECT 17.990 171.715 18.270 171.750 ;
        RECT 31.580 166.650 31.880 171.800 ;
        RECT 35.730 169.300 38.010 169.600 ;
        RECT 35.730 168.600 36.030 169.300 ;
        RECT 35.730 168.300 42.660 168.600 ;
        RECT 19.090 166.500 19.370 166.535 ;
        RECT 19.080 166.200 26.010 166.500 ;
        RECT 31.580 166.350 33.960 166.650 ;
        RECT 19.090 166.165 19.370 166.200 ;
        RECT 21.030 164.300 21.330 166.200 ;
        RECT 31.580 164.300 31.880 166.350 ;
        RECT 35.730 164.300 36.030 168.300 ;
        RECT 21.030 164.000 36.030 164.300 ;
        RECT 21.030 157.850 21.330 164.000 ;
        RECT 35.730 161.000 36.030 164.000 ;
        RECT 35.730 160.700 49.110 161.000 ;
        RECT 35.730 158.250 36.030 160.700 ;
        RECT 47.230 160.050 47.530 160.700 ;
        RECT 47.230 159.750 55.960 160.050 ;
        RECT 33.600 157.950 36.030 158.250 ;
        RECT 21.030 157.550 25.910 157.850 ;
        RECT 21.030 153.100 21.330 157.550 ;
        RECT 35.730 155.950 36.030 157.950 ;
        RECT 35.730 155.650 38.610 155.950 ;
        RECT 37.430 155.050 37.730 155.650 ;
        RECT 43.050 155.050 43.415 155.055 ;
        RECT 37.430 154.750 43.415 155.050 ;
        RECT 21.030 152.800 29.910 153.100 ;
        RECT 21.030 141.750 21.330 152.800 ;
        RECT 28.730 151.750 29.030 152.800 ;
        RECT 32.630 151.750 32.930 152.630 ;
        RECT 28.730 151.450 32.930 151.750 ;
        RECT 31.130 142.250 36.210 142.550 ;
        RECT 31.130 142.050 31.430 142.250 ;
        RECT 28.450 141.750 31.430 142.050 ;
        RECT 21.030 141.450 23.460 141.750 ;
        RECT 21.030 139.500 21.330 141.450 ;
        RECT 31.130 140.450 31.430 141.750 ;
        RECT 39.980 140.450 40.280 141.730 ;
        RECT 31.130 140.150 50.560 140.450 ;
        RECT 31.130 139.500 31.430 140.150 ;
        RECT 21.030 139.200 31.430 139.500 ;
        RECT 49.530 138.950 49.830 140.150 ;
        RECT 54.830 139.450 56.310 139.750 ;
        RECT 54.830 138.950 55.130 139.450 ;
        RECT 49.530 138.650 55.130 138.950 ;
      LAYER met3 ;
        RECT 17.965 172.050 18.295 172.065 ;
        RECT 9.580 171.750 18.295 172.050 ;
        RECT 9.580 168.150 9.880 171.750 ;
        RECT 17.965 171.735 18.295 171.750 ;
        RECT 9.580 167.850 13.080 168.150 ;
        RECT 3.000 166.500 5.060 167.350 ;
        RECT 12.780 166.500 13.080 167.850 ;
        RECT 19.065 166.500 19.395 166.515 ;
        RECT 3.000 166.200 19.395 166.500 ;
        RECT 3.000 165.350 5.060 166.200 ;
        RECT 19.065 166.185 19.395 166.200 ;
      LAYER met4 ;
        RECT 3.030 167.355 5.030 220.760 ;
        RECT 3.025 165.345 5.035 167.355 ;
        RECT 3.030 5.000 5.030 165.345 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 30.940 172.655 31.870 173.565 ;
        RECT 30.940 172.635 31.045 172.655 ;
        RECT 30.875 172.465 31.045 172.635 ;
        RECT 38.335 169.655 39.685 170.565 ;
        RECT 38.480 169.465 38.650 169.655 ;
        RECT 30.490 167.355 31.420 168.265 ;
        RECT 30.490 167.335 30.595 167.355 ;
        RECT 30.425 167.165 30.595 167.335 ;
        RECT 49.765 161.045 52.935 161.955 ;
        RECT 49.865 160.855 50.035 161.045 ;
        RECT 29.440 158.505 30.370 159.415 ;
        RECT 29.440 158.485 29.545 158.505 ;
        RECT 29.375 158.315 29.545 158.485 ;
        RECT 39.085 156.005 40.435 156.915 ;
        RECT 39.230 155.815 39.400 156.005 ;
        RECT 29.480 153.645 30.410 154.555 ;
        RECT 29.480 153.625 29.585 153.645 ;
        RECT 29.415 153.455 29.585 153.625 ;
        RECT 22.870 143.035 24.675 143.265 ;
        RECT 22.385 142.355 24.675 143.035 ;
        RECT 36.880 142.595 37.810 143.505 ;
        RECT 36.880 142.575 36.985 142.595 ;
        RECT 36.815 142.405 36.985 142.575 ;
        RECT 22.530 142.165 22.700 142.355 ;
        RECT 51.420 141.185 53.225 141.415 ;
        RECT 50.935 140.505 53.225 141.185 ;
        RECT 51.080 140.315 51.250 140.505 ;
      LAYER li1 ;
        RECT 31.450 174.035 31.780 175.015 ;
        RECT 31.550 173.715 31.780 174.035 ;
        RECT 31.550 173.485 33.145 173.715 ;
        RECT 31.550 173.435 31.780 173.485 ;
        RECT 31.450 172.805 31.780 173.435 ;
        RECT 37.680 172.900 38.330 173.100 ;
        RECT 37.680 171.750 37.880 172.900 ;
        RECT 38.425 171.750 38.755 172.000 ;
        RECT 37.680 171.550 38.755 171.750 ;
        RECT 38.425 171.215 38.755 171.550 ;
        RECT 38.425 171.045 39.105 171.215 ;
        RECT 38.415 170.625 38.765 170.875 ;
        RECT 38.935 170.445 39.105 171.045 ;
        RECT 39.275 170.845 39.625 170.875 ;
        RECT 39.275 170.655 40.825 170.845 ;
        RECT 39.275 170.625 39.625 170.655 ;
        RECT 38.845 169.805 39.175 170.445 ;
        RECT 31.000 168.735 31.330 169.715 ;
        RECT 30.600 168.550 30.930 168.565 ;
        RECT 29.480 168.350 30.930 168.550 ;
        RECT 30.600 168.325 30.930 168.350 ;
        RECT 31.100 168.415 31.330 168.735 ;
        RECT 31.100 168.185 32.595 168.415 ;
        RECT 31.100 168.135 31.330 168.185 ;
        RECT 31.000 167.505 31.330 168.135 ;
        RECT 49.805 162.725 50.185 163.405 ;
        RECT 51.115 162.895 51.445 163.405 ;
        RECT 51.955 162.895 52.355 163.405 ;
        RECT 51.115 162.725 52.355 162.895 ;
        RECT 52.535 162.750 52.855 163.405 ;
        RECT 49.805 161.765 49.975 162.725 ;
        RECT 50.145 162.385 51.450 162.555 ;
        RECT 52.535 162.475 52.930 162.750 ;
        RECT 50.145 161.935 50.390 162.385 ;
        RECT 50.560 162.015 51.110 162.215 ;
        RECT 51.280 162.185 51.450 162.385 ;
        RECT 52.225 162.450 52.930 162.475 ;
        RECT 52.225 162.305 52.855 162.450 ;
        RECT 51.280 162.015 51.655 162.185 ;
        RECT 51.825 161.765 52.055 162.265 ;
        RECT 49.805 161.595 52.055 161.765 ;
        RECT 50.355 161.275 50.525 161.595 ;
        RECT 52.225 161.425 52.395 162.305 ;
        RECT 51.440 161.255 52.395 161.425 ;
        RECT 29.950 159.885 30.280 160.865 ;
        RECT 30.050 159.515 30.280 159.885 ;
        RECT 30.050 159.285 31.595 159.515 ;
        RECT 29.950 158.655 30.280 159.285 ;
        RECT 31.365 159.135 31.595 159.285 ;
        RECT 39.175 158.100 39.505 158.350 ;
        RECT 39.030 157.800 39.505 158.100 ;
        RECT 39.175 157.565 39.505 157.800 ;
        RECT 39.175 157.395 39.855 157.565 ;
        RECT 38.105 156.975 39.515 157.225 ;
        RECT 39.685 156.795 39.855 157.395 ;
        RECT 40.025 157.200 40.375 157.225 ;
        RECT 40.025 157.000 41.330 157.200 ;
        RECT 40.025 156.975 40.375 157.000 ;
        RECT 39.595 156.155 39.925 156.795 ;
        RECT 29.990 155.025 30.320 156.005 ;
        RECT 29.590 154.850 29.920 154.855 ;
        RECT 28.430 154.650 29.920 154.850 ;
        RECT 29.590 154.615 29.920 154.650 ;
        RECT 30.090 154.665 30.320 155.025 ;
        RECT 31.365 154.665 31.595 154.915 ;
        RECT 30.090 154.435 31.595 154.665 ;
        RECT 30.090 154.425 30.320 154.435 ;
        RECT 29.990 153.795 30.320 154.425 ;
        RECT 22.465 144.315 22.725 144.715 ;
        RECT 24.000 144.375 24.595 144.715 ;
        RECT 22.465 144.145 23.830 144.315 ;
        RECT 22.465 143.500 22.925 143.975 ;
        RECT 21.630 143.300 22.925 143.500 ;
        RECT 22.465 143.245 22.925 143.300 ;
        RECT 23.095 143.075 23.830 144.145 ;
        RECT 22.465 142.905 23.830 143.075 ;
        RECT 24.000 143.055 24.175 144.375 ;
        RECT 24.355 143.450 24.595 144.205 ;
        RECT 37.390 143.975 37.720 144.955 ;
        RECT 36.990 143.800 37.320 143.805 ;
        RECT 35.880 143.600 37.320 143.800 ;
        RECT 36.990 143.565 37.320 143.600 ;
        RECT 24.355 143.250 25.530 143.450 ;
        RECT 37.490 143.375 37.720 143.975 ;
        RECT 24.355 143.225 24.595 143.250 ;
        RECT 22.465 142.505 22.725 142.905 ;
        RECT 24.000 142.505 24.595 143.055 ;
        RECT 37.390 142.745 37.720 143.375 ;
        RECT 51.015 142.465 51.275 142.865 ;
        RECT 51.015 142.295 52.380 142.465 ;
        RECT 51.015 141.650 51.475 142.125 ;
        RECT 50.130 141.450 51.475 141.650 ;
        RECT 51.015 141.395 51.475 141.450 ;
        RECT 51.645 141.225 52.380 142.295 ;
        RECT 52.905 141.650 53.145 142.355 ;
        RECT 52.905 141.450 54.230 141.650 ;
        RECT 52.905 141.375 53.145 141.450 ;
        RECT 51.015 141.055 52.380 141.225 ;
        RECT 51.015 140.655 51.275 141.055 ;
      LAYER met1 ;
        RECT 149.100 225.450 161.000 225.750 ;
        RECT 149.100 225.400 149.400 225.450 ;
        RECT 32.915 178.285 37.395 178.515 ;
        RECT 32.915 173.455 33.145 178.285 ;
        RECT 32.365 171.185 36.395 171.415 ;
        RECT 29.435 168.550 29.725 168.565 ;
        RECT 24.480 168.350 29.725 168.550 ;
        RECT 24.480 154.850 24.680 168.350 ;
        RECT 29.435 168.335 29.725 168.350 ;
        RECT 32.365 168.155 32.595 171.185 ;
        RECT 36.165 168.665 36.395 171.185 ;
        RECT 37.165 170.865 37.395 178.285 ;
        RECT 40.080 173.900 44.630 174.100 ;
        RECT 38.035 173.100 38.325 173.115 ;
        RECT 40.080 173.100 40.280 173.900 ;
        RECT 38.030 172.900 40.280 173.100 ;
        RECT 38.035 172.885 38.325 172.900 ;
        RECT 37.165 170.635 38.775 170.865 ;
        RECT 40.615 168.665 40.845 170.895 ;
        RECT 36.165 168.435 40.845 168.665 ;
        RECT 31.365 162.535 37.695 162.765 ;
        RECT 31.365 159.155 31.595 162.535 ;
        RECT 31.365 157.285 35.845 157.515 ;
        RECT 28.385 154.850 28.675 154.865 ;
        RECT 24.480 154.650 28.675 154.850 ;
        RECT 31.365 154.820 31.595 157.285 ;
        RECT 24.480 149.000 24.680 154.650 ;
        RECT 28.385 154.635 28.675 154.650 ;
        RECT 31.360 154.580 31.600 154.820 ;
        RECT 31.365 154.435 31.595 154.580 ;
        RECT 35.615 154.515 35.845 157.285 ;
        RECT 37.465 157.215 37.695 162.535 ;
        RECT 44.430 162.550 44.630 173.900 ;
        RECT 47.230 166.350 60.080 166.550 ;
        RECT 47.230 162.550 47.430 166.350 ;
        RECT 52.580 162.550 54.330 162.750 ;
        RECT 44.430 162.350 49.080 162.550 ;
        RECT 52.610 162.470 52.930 162.550 ;
        RECT 48.805 162.335 49.080 162.350 ;
        RECT 48.805 162.275 50.305 162.335 ;
        RECT 48.805 162.185 50.375 162.275 ;
        RECT 50.085 162.045 50.375 162.185 ;
        RECT 50.530 162.200 50.760 162.275 ;
        RECT 50.530 162.050 51.105 162.200 ;
        RECT 50.530 161.985 50.760 162.050 ;
        RECT 50.530 161.700 50.730 161.985 ;
        RECT 38.280 161.500 50.730 161.700 ;
        RECT 38.280 158.050 38.480 161.500 ;
        RECT 39.085 158.050 39.345 158.080 ;
        RECT 38.280 157.850 39.430 158.050 ;
        RECT 39.085 157.820 39.345 157.850 ;
        RECT 38.225 157.215 38.535 157.225 ;
        RECT 37.465 156.985 38.535 157.215 ;
        RECT 41.035 156.985 41.995 157.215 ;
        RECT 38.225 156.975 38.535 156.985 ;
        RECT 41.765 154.515 41.995 156.985 ;
        RECT 35.615 154.285 41.995 154.515 ;
        RECT 54.130 150.500 54.330 162.550 ;
        RECT 19.130 148.800 24.680 149.000 ;
        RECT 35.880 150.300 54.330 150.500 ;
        RECT 19.130 140.100 19.330 148.800 ;
        RECT 21.630 146.550 34.180 146.750 ;
        RECT 21.630 143.545 21.830 146.550 ;
        RECT 21.615 143.255 21.845 143.545 ;
        RECT 25.285 143.450 25.575 143.465 ;
        RECT 25.285 143.250 26.780 143.450 ;
        RECT 25.285 143.235 25.575 143.250 ;
        RECT 24.335 142.900 24.625 142.915 ;
        RECT 24.335 142.700 25.830 142.900 ;
        RECT 24.335 142.685 24.625 142.700 ;
        RECT 25.630 140.100 25.830 142.700 ;
        RECT 26.580 141.300 26.780 143.250 ;
        RECT 26.580 141.100 31.430 141.300 ;
        RECT 19.130 139.900 25.830 140.100 ;
        RECT 31.230 139.050 31.430 141.100 ;
        RECT 33.980 141.150 34.180 146.550 ;
        RECT 35.880 143.860 36.080 150.300 ;
        RECT 35.850 143.540 36.110 143.860 ;
        RECT 37.435 143.700 37.725 143.715 ;
        RECT 37.435 143.500 39.380 143.700 ;
        RECT 37.435 143.485 37.725 143.500 ;
        RECT 39.180 141.150 39.380 143.500 ;
        RECT 42.680 142.150 42.880 150.300 ;
        RECT 59.880 148.550 60.080 166.350 ;
        RECT 45.430 148.350 60.080 148.550 ;
        RECT 45.430 145.050 45.630 148.350 ;
        RECT 45.430 144.850 54.230 145.050 ;
        RECT 44.350 142.150 44.610 142.210 ;
        RECT 42.680 141.950 44.610 142.150 ;
        RECT 44.350 141.890 44.610 141.950 ;
        RECT 33.980 140.950 39.380 141.150 ;
        RECT 45.430 139.050 45.630 144.850 ;
        RECT 46.450 142.150 46.710 142.210 ;
        RECT 46.450 141.950 50.330 142.150 ;
        RECT 46.450 141.890 46.710 141.950 ;
        RECT 50.130 141.695 50.330 141.950 ;
        RECT 54.030 141.695 54.230 144.850 ;
        RECT 50.115 141.405 50.345 141.695 ;
        RECT 54.015 141.405 54.245 141.695 ;
        RECT 31.230 138.850 45.630 139.050 ;
      LAYER met2 ;
        RECT 44.320 142.150 44.640 142.180 ;
        RECT 46.420 142.150 46.740 142.180 ;
        RECT 44.320 141.950 46.740 142.150 ;
        RECT 44.320 141.920 44.640 141.950 ;
        RECT 46.420 141.920 46.740 141.950 ;
  END
END tt_um_test_17
END LIBRARY

