VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_template
  CLASS BLOCK ;
  FOREIGN tt_um_template ;
  ORIGIN 0.000 0.000 ;
  SIZE 151.710 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 142.830 224.760 143.130 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 142.975 225.255 142.985 225.265 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 145.590 224.760 145.890 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.735 225.255 145.745 225.265 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 140.070 224.760 140.370 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.215 225.255 140.225 225.265 ;
    END
  END rst_n
  PIN ua[0]
    PORT
      LAYER met4 ;
        RECT 150.810 0.000 151.710 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.255 0.495 151.265 0.505 ;
    END
  END ua[0]
  PIN ua[1]
    PORT
      LAYER met4 ;
        RECT 131.490 0.000 132.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT 112.170 0.000 113.070 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.615 0.495 112.625 0.505 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 92.850 0.000 93.750 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.295 0.495 93.305 0.505 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 73.530 0.000 74.430 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.975 0.495 73.985 0.505 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 54.210 0.000 55.110 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.655 0.495 54.665 0.505 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 34.890 0.000 35.790 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.335 0.495 35.345 0.505 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 15.570 0.000 16.470 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.015 0.495 16.025 0.505 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 137.310 224.760 137.610 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.455 225.255 137.465 225.265 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 134.550 224.760 134.850 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.695 225.255 134.705 225.265 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 131.790 224.760 132.090 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.935 225.255 131.945 225.265 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 129.030 224.760 129.330 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.175 225.255 129.185 225.265 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 126.270 224.760 126.570 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.415 225.255 126.425 225.265 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 123.510 224.760 123.810 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.655 225.255 123.665 225.265 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 120.750 224.760 121.050 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.895 225.255 120.905 225.265 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 117.990 224.760 118.290 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.135 225.255 118.145 225.265 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 115.230 224.760 115.530 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.375 225.255 115.385 225.265 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 112.470 224.760 112.770 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.615 225.255 112.625 225.265 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 109.710 224.760 110.010 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.855 225.255 109.865 225.265 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 106.950 224.760 107.250 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.095 225.255 107.105 225.265 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 104.190 224.760 104.490 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.335 225.255 104.345 225.265 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 101.430 224.760 101.730 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.575 225.255 101.585 225.265 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 98.670 224.760 98.970 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.815 225.255 98.825 225.265 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 95.910 224.760 96.210 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.055 225.255 96.065 225.265 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 48.990 224.760 49.290 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.135 225.255 49.145 225.265 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 46.230 224.760 46.530 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.375 225.255 46.385 225.265 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 43.470 224.760 43.770 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.615 225.255 43.625 225.265 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 40.710 224.760 41.010 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.855 225.255 40.865 225.265 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 37.950 224.760 38.250 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.095 225.255 38.105 225.265 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 35.190 224.760 35.490 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.335 225.255 35.345 225.265 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 32.430 224.760 32.730 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.575 225.255 32.585 225.265 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 29.670 224.760 29.970 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.815 225.255 29.825 225.265 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 71.070 224.760 71.370 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.215 225.255 71.225 225.265 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 68.310 224.760 68.610 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.455 225.255 68.465 225.265 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 65.550 224.760 65.850 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.695 225.255 65.705 225.265 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 62.790 224.760 63.090 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.935 225.255 62.945 225.265 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 60.030 224.760 60.330 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.175 225.255 60.185 225.265 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 57.270 224.760 57.570 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.415 225.255 57.425 225.265 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 54.510 224.760 54.810 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.655 225.255 54.665 225.265 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 51.750 224.760 52.050 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.895 225.255 51.905 225.265 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 93.150 224.760 93.450 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.295 225.255 93.305 225.265 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 90.390 224.760 90.690 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.535 225.255 90.545 225.265 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 87.630 224.760 87.930 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.775 225.255 87.785 225.265 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 84.870 224.760 85.170 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.015 225.255 85.025 225.265 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 82.110 224.760 82.410 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.255 225.255 82.265 225.265 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 79.350 224.760 79.650 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.495 225.255 79.505 225.265 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 76.590 224.760 76.890 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.735 225.255 76.745 225.265 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 73.830 224.760 74.130 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.975 225.255 73.985 225.265 ;
    END
  END uo_out[7]
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 0.000 5.000 2.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.000 5.000 5.000 220.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 22.440 189.105 57.650 215.905 ;
      LAYER met1 ;
        RECT 7.145 187.265 65.725 218.580 ;
      LAYER met2 ;
        RECT 6.030 6.920 151.475 218.625 ;
      LAYER met3 ;
        RECT 1.610 0.130 151.590 218.645 ;
      LAYER met4 ;
        RECT 2.400 206.980 2.600 218.550 ;
        RECT 5.400 206.980 6.895 218.550 ;
  END
END tt_um_template
END LIBRARY

