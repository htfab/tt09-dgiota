VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_5
  CLASS BLOCK ;
  FOREIGN tt_um_test_5 ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.510 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 142.830 224.760 143.130 225.760 ;
    END
  END clk
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2.445 131.235 2.755 131.305 ;
        RECT 1.340 131.210 2.810 131.235 ;
        RECT 1.340 130.885 2.860 131.210 ;
        RECT 1.340 130.515 2.810 130.885 ;
        RECT 2.175 130.220 2.725 130.515 ;
        RECT 2.175 130.070 2.580 130.220 ;
      LAYER via3 ;
        RECT 1.400 130.625 1.900 131.125 ;
      LAYER met4 ;
        RECT 0.000 5.000 2.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.590 224.760 145.890 225.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3.350 134.815 5.350 135.630 ;
        RECT 9.975 134.815 10.675 134.825 ;
        RECT 3.350 134.625 10.675 134.815 ;
        RECT 3.350 134.385 10.925 134.625 ;
        RECT 3.350 133.570 5.350 134.385 ;
        RECT 10.375 134.325 10.925 134.385 ;
        RECT 10.375 134.320 10.875 134.325 ;
        RECT 10.375 134.125 10.825 134.320 ;
      LAYER via3 ;
        RECT 3.350 133.600 5.350 135.600 ;
      LAYER met4 ;
        RECT 3.000 135.605 5.000 220.760 ;
        RECT 3.000 133.595 5.355 135.605 ;
        RECT 3.000 5.000 5.000 133.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.070 224.760 140.370 225.760 ;
    END
  END VGND
  PIN ua[0]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.471000 ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER li1 ;
        RECT 68.855 154.745 69.175 155.455 ;
        RECT 68.855 154.560 71.140 154.745 ;
        RECT 68.855 154.525 69.175 154.560 ;
        RECT 68.545 154.355 69.175 154.525 ;
        RECT 68.545 153.475 68.715 154.355 ;
        RECT 67.760 153.305 68.715 153.475 ;
        RECT 49.770 140.015 51.335 140.185 ;
        RECT 49.770 139.945 50.100 140.015 ;
        RECT 68.485 135.790 68.945 136.225 ;
        RECT 68.160 135.605 68.945 135.790 ;
        RECT 68.485 135.495 68.945 135.605 ;
      LAYER mcon ;
        RECT 70.955 154.560 71.140 154.745 ;
        RECT 51.165 140.015 51.335 140.185 ;
        RECT 68.170 135.615 68.340 135.785 ;
      LAYER met1 ;
        RECT 70.925 154.685 71.170 154.805 ;
        RECT 72.470 154.685 72.730 154.760 ;
        RECT 70.925 154.515 72.785 154.685 ;
        RECT 70.925 154.500 71.170 154.515 ;
        RECT 51.105 139.985 51.395 140.215 ;
        RECT 51.165 136.495 51.335 139.985 ;
        RECT 70.955 138.145 71.140 154.500 ;
        RECT 72.470 154.440 72.730 154.515 ;
        RECT 54.210 137.960 71.140 138.145 ;
        RECT 54.210 136.495 54.395 137.960 ;
        RECT 51.160 136.310 54.395 136.495 ;
        RECT 66.060 135.790 66.245 137.960 ;
        RECT 68.110 135.790 68.400 135.815 ;
        RECT 66.060 135.605 68.400 135.790 ;
        RECT 68.110 135.585 68.400 135.605 ;
      LAYER via ;
        RECT 72.470 154.470 72.730 154.730 ;
      LAYER met2 ;
        RECT 72.440 154.685 72.760 154.730 ;
        RECT 72.440 154.515 149.085 154.685 ;
        RECT 72.440 154.470 72.760 154.515 ;
        RECT 148.915 5.285 149.085 154.515 ;
        RECT 150.395 5.285 150.805 5.310 ;
        RECT 148.915 5.115 150.805 5.285 ;
        RECT 150.395 5.030 150.805 5.115 ;
      LAYER via2 ;
        RECT 150.440 5.030 150.760 5.310 ;
      LAYER met3 ;
        RECT 150.415 4.965 151.785 5.335 ;
        RECT 151.415 3.385 151.785 4.965 ;
        RECT 151.115 3.015 151.785 3.385 ;
        RECT 151.115 2.315 151.485 3.015 ;
      LAYER via3 ;
        RECT 151.115 2.365 151.485 2.735 ;
      LAYER met4 ;
        RECT 151.110 2.360 151.490 2.740 ;
        RECT 151.115 1.000 151.485 2.360 ;
        RECT 150.810 0.000 151.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 51.820 158.640 52.150 158.665 ;
        RECT 51.565 158.465 52.150 158.640 ;
        RECT 51.820 158.425 52.150 158.465 ;
      LAYER mcon ;
        RECT 51.615 158.470 51.785 158.640 ;
      LAYER met1 ;
        RECT 51.045 158.640 51.365 158.685 ;
        RECT 51.555 158.640 51.845 158.670 ;
        RECT 51.045 158.465 51.845 158.640 ;
        RECT 51.045 158.425 51.365 158.465 ;
        RECT 51.555 158.440 51.845 158.465 ;
      LAYER via ;
        RECT 51.075 158.425 51.335 158.685 ;
      LAYER met2 ;
        RECT 34.715 169.110 160.385 169.285 ;
        RECT 34.715 158.640 34.890 169.110 ;
        RECT 51.075 158.640 51.335 158.715 ;
        RECT 34.715 158.465 51.340 158.640 ;
        RECT 51.075 158.395 51.335 158.465 ;
        RECT 160.210 127.465 160.385 169.110 ;
        RECT 160.085 127.185 160.510 127.465 ;
        RECT 160.210 127.145 160.385 127.185 ;
      LAYER via2 ;
        RECT 160.130 127.185 160.465 127.465 ;
      LAYER met3 ;
        RECT 160.105 40.655 160.490 127.490 ;
        RECT 131.760 40.270 160.490 40.655 ;
        RECT 131.760 1.785 132.145 40.270 ;
        RECT 131.755 1.325 132.155 1.785 ;
      LAYER via3 ;
        RECT 131.755 1.355 132.155 1.755 ;
      LAYER met4 ;
        RECT 131.835 1.760 132.235 1.870 ;
        RECT 131.750 1.435 132.235 1.760 ;
        RECT 131.750 1.350 132.270 1.435 ;
        RECT 131.835 1.000 132.270 1.350 ;
        RECT 131.490 0.000 132.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 65.920 144.365 66.250 144.385 ;
        RECT 65.920 144.155 67.005 144.365 ;
        RECT 65.920 144.145 66.250 144.155 ;
      LAYER mcon ;
        RECT 66.795 144.155 67.005 144.365 ;
      LAYER met1 ;
        RECT 66.765 144.365 67.035 144.425 ;
        RECT 69.970 144.365 70.230 144.420 ;
        RECT 66.745 144.155 70.230 144.365 ;
        RECT 66.765 144.095 67.035 144.155 ;
        RECT 69.970 144.100 70.230 144.155 ;
      LAYER via ;
        RECT 69.970 144.130 70.230 144.390 ;
      LAYER met2 ;
        RECT 69.940 144.365 70.260 144.390 ;
        RECT 69.940 144.155 111.205 144.365 ;
        RECT 69.940 144.130 70.260 144.155 ;
        RECT 110.995 5.375 111.205 144.155 ;
        RECT 110.880 5.095 111.320 5.375 ;
        RECT 110.995 4.745 111.205 5.095 ;
      LAYER via2 ;
        RECT 110.925 5.095 111.275 5.375 ;
      LAYER met3 ;
        RECT 110.900 4.700 111.300 5.400 ;
        RECT 110.900 4.300 112.900 4.700 ;
        RECT 112.500 2.400 112.900 4.300 ;
      LAYER via3 ;
        RECT 112.500 2.450 112.900 2.850 ;
      LAYER met4 ;
        RECT 112.495 2.445 112.905 2.855 ;
        RECT 112.500 1.000 112.900 2.445 ;
        RECT 112.170 0.000 113.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 92.850 0.000 93.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 73.530 0.000 74.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 54.210 0.000 55.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 34.890 0.000 35.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 15.570 0.000 16.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 137.310 224.760 137.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 134.550 224.760 134.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 131.790 224.760 132.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 129.030 224.760 129.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 126.270 224.760 126.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 123.510 224.760 123.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 120.750 224.760 121.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 117.990 224.760 118.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 115.230 224.760 115.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 112.470 224.760 112.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 109.710 224.760 110.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 106.950 224.760 107.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 104.190 224.760 104.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 101.430 224.760 101.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 98.670 224.760 98.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 95.910 224.760 96.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 48.990 224.760 49.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 46.230 224.760 46.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 43.470 224.760 43.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 40.710 224.760 41.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 37.950 224.760 38.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 35.190 224.760 35.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 32.430 224.760 32.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 29.670 224.760 29.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 71.070 224.760 71.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 68.310 224.760 68.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 65.550 224.760 65.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 62.790 224.760 63.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 60.030 224.760 60.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 57.270 224.760 57.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 54.510 224.760 54.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 51.750 224.760 52.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 93.150 224.760 93.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 90.390 224.760 90.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 87.630 224.760 87.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 84.870 224.760 85.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 82.110 224.760 82.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 79.350 224.760 79.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 76.590 224.760 76.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 73.830 224.760 74.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 53.385 160.765 53.555 161.290 ;
      LAYER nwell ;
        RECT 53.050 160.260 53.890 160.305 ;
        RECT 51.310 158.700 53.890 160.260 ;
      LAYER pwell ;
        RECT 57.485 159.165 57.655 159.690 ;
      LAYER nwell ;
        RECT 51.310 158.655 53.070 158.700 ;
        RECT 57.150 158.500 57.990 158.705 ;
      LAYER pwell ;
        RECT 51.645 157.265 51.815 157.435 ;
      LAYER nwell ;
        RECT 57.150 157.100 59.660 158.500 ;
      LAYER pwell ;
        RECT 69.735 157.115 69.905 157.640 ;
      LAYER nwell ;
        RECT 57.900 156.895 59.660 157.100 ;
        RECT 69.400 155.900 70.240 156.655 ;
      LAYER pwell ;
        RECT 59.150 155.505 59.320 155.675 ;
      LAYER nwell ;
        RECT 65.850 155.050 70.240 155.900 ;
        RECT 65.850 154.295 69.450 155.050 ;
      LAYER pwell ;
        RECT 66.185 152.905 66.355 153.075 ;
      LAYER nwell ;
        RECT 59.360 150.340 60.965 152.020 ;
      LAYER pwell ;
        RECT 62.185 150.595 62.355 150.765 ;
      LAYER nwell ;
        RECT 58.795 150.260 60.965 150.340 ;
      LAYER pwell ;
        RECT 57.810 149.835 58.335 150.005 ;
      LAYER nwell ;
        RECT 58.795 149.500 60.400 150.260 ;
      LAYER pwell ;
        RECT 60.235 147.715 60.405 148.240 ;
        RECT 52.685 146.665 52.855 147.190 ;
      LAYER nwell ;
        RECT 52.350 146.150 53.190 146.205 ;
        RECT 52.350 144.600 54.760 146.150 ;
        RECT 59.900 145.650 60.740 147.255 ;
        RECT 53.000 144.545 54.760 144.600 ;
        RECT 59.050 144.045 60.810 145.650 ;
      LAYER pwell ;
        RECT 66.255 145.375 66.425 145.545 ;
      LAYER nwell ;
        RECT 65.000 143.550 66.760 144.155 ;
      LAYER pwell ;
        RECT 53.335 143.155 53.505 143.325 ;
        RECT 59.390 142.655 59.560 142.825 ;
      LAYER nwell ;
        RECT 65.000 142.550 67.490 143.550 ;
        RECT 66.650 141.945 67.490 142.550 ;
      LAYER pwell ;
        RECT 50.105 141.175 50.275 141.345 ;
        RECT 66.985 140.960 67.155 141.485 ;
      LAYER nwell ;
        RECT 48.850 139.300 50.610 139.955 ;
        RECT 48.850 138.350 51.190 139.300 ;
        RECT 50.350 137.695 51.190 138.350 ;
      LAYER pwell ;
        RECT 50.685 136.710 50.855 137.235 ;
      LAYER nwell ;
        RECT 68.210 136.940 70.890 137.410 ;
      LAYER pwell ;
        RECT 46.380 136.525 46.550 136.695 ;
      LAYER nwell ;
        RECT 68.210 136.100 72.455 136.940 ;
      LAYER pwell ;
        RECT 72.915 136.435 73.440 136.605 ;
      LAYER nwell ;
        RECT 68.210 135.805 70.890 136.100 ;
        RECT 44.210 134.650 46.890 135.305 ;
        RECT 44.210 133.810 48.495 134.650 ;
      LAYER pwell ;
        RECT 68.550 134.415 68.720 134.585 ;
        RECT 48.955 134.145 49.480 134.315 ;
      LAYER nwell ;
        RECT 44.210 133.700 46.890 133.810 ;
      LAYER li1 ;
        RECT 53.240 161.525 53.700 161.695 ;
        RECT 53.325 160.800 53.615 161.525 ;
        RECT 51.500 159.985 52.880 160.155 ;
        RECT 51.840 158.845 52.050 159.985 ;
        RECT 52.220 158.835 52.550 159.815 ;
        RECT 53.325 158.975 53.615 160.140 ;
        RECT 57.340 159.925 57.800 160.095 ;
        RECT 57.425 159.200 57.715 159.925 ;
        RECT 52.320 158.495 52.550 158.835 ;
        RECT 53.240 158.805 53.700 158.975 ;
        RECT 52.880 158.495 54.085 158.590 ;
        RECT 52.320 158.415 54.085 158.495 ;
        RECT 52.320 158.310 53.040 158.415 ;
        RECT 51.820 157.435 52.050 158.255 ;
        RECT 52.320 158.235 52.550 158.310 ;
        RECT 52.220 157.605 52.550 158.235 ;
        RECT 53.910 157.585 54.085 158.415 ;
        RECT 51.500 157.265 52.880 157.435 ;
        RECT 53.910 157.415 54.090 157.585 ;
        RECT 53.910 157.090 54.085 157.415 ;
        RECT 57.425 157.375 57.715 158.540 ;
        RECT 58.090 158.225 59.470 158.395 ;
        RECT 57.340 157.205 57.800 157.375 ;
        RECT 55.910 156.845 56.095 157.090 ;
        RECT 58.185 157.085 58.515 158.225 ;
        RECT 59.045 157.255 59.375 158.040 ;
        RECT 69.590 157.875 70.050 158.045 ;
        RECT 58.695 157.085 59.375 157.255 ;
        RECT 69.675 157.150 69.965 157.875 ;
        RECT 58.175 156.845 58.525 156.915 ;
        RECT 55.910 156.665 58.525 156.845 ;
        RECT 55.910 156.660 58.320 156.665 ;
        RECT 58.695 156.485 58.865 157.085 ;
        RECT 59.035 156.840 59.385 156.915 ;
        RECT 59.035 156.665 59.640 156.840 ;
        RECT 59.245 156.660 59.640 156.665 ;
        RECT 58.185 155.675 58.455 156.485 ;
        RECT 58.625 155.845 58.955 156.485 ;
        RECT 59.125 155.675 59.365 156.485 ;
        RECT 58.090 155.505 59.470 155.675 ;
        RECT 66.040 155.625 69.260 155.795 ;
        RECT 66.125 154.775 66.505 155.455 ;
        RECT 66.125 153.815 66.295 154.775 ;
        RECT 66.715 154.605 66.885 155.035 ;
        RECT 67.095 154.775 67.265 155.625 ;
        RECT 67.435 154.945 67.765 155.455 ;
        RECT 67.935 155.115 68.105 155.625 ;
        RECT 68.275 154.945 68.675 155.455 ;
        RECT 69.675 155.325 69.965 156.490 ;
        RECT 69.590 155.155 70.050 155.325 ;
        RECT 67.435 154.775 68.675 154.945 ;
        RECT 66.465 154.435 67.770 154.605 ;
        RECT 66.465 153.985 66.710 154.435 ;
        RECT 66.880 154.065 67.430 154.265 ;
        RECT 67.600 154.235 67.770 154.435 ;
        RECT 67.600 154.065 67.975 154.235 ;
        RECT 68.145 153.815 68.375 154.315 ;
        RECT 66.125 153.645 68.375 153.815 ;
        RECT 66.175 153.075 66.505 153.465 ;
        RECT 66.675 153.325 66.845 153.645 ;
        RECT 67.015 153.075 67.345 153.465 ;
        RECT 68.885 153.075 69.175 153.910 ;
        RECT 66.040 152.905 69.260 153.075 ;
        RECT 59.465 151.000 59.635 151.830 ;
        RECT 61.365 151.500 61.635 151.595 ;
        RECT 59.805 151.270 62.015 151.500 ;
        RECT 59.805 151.170 60.785 151.270 ;
        RECT 61.385 151.170 62.015 151.270 ;
        RECT 59.465 150.790 60.775 151.000 ;
        RECT 59.465 150.450 59.635 150.790 ;
        RECT 60.955 150.770 61.195 151.100 ;
        RECT 62.185 151.000 62.355 151.830 ;
        RECT 61.365 150.770 62.355 151.000 ;
        RECT 62.185 150.450 62.355 150.770 ;
        RECT 57.405 150.065 57.575 150.150 ;
        RECT 60.125 150.065 60.295 150.150 ;
        RECT 57.405 149.775 58.300 150.065 ;
        RECT 58.960 149.775 60.295 150.065 ;
        RECT 57.405 149.690 57.575 149.775 ;
        RECT 60.125 149.690 60.295 149.775 ;
        RECT 60.090 148.475 60.550 148.645 ;
        RECT 60.175 147.750 60.465 148.475 ;
        RECT 52.540 147.425 53.000 147.595 ;
        RECT 52.625 146.700 52.915 147.425 ;
        RECT 55.385 146.480 55.610 146.610 ;
        RECT 55.790 146.480 58.270 146.490 ;
        RECT 55.385 146.255 58.270 146.480 ;
        RECT 52.625 144.875 52.915 146.040 ;
        RECT 53.190 145.875 54.570 146.045 ;
        RECT 53.275 144.905 53.535 145.875 ;
        RECT 52.540 144.705 53.000 144.875 ;
        RECT 53.275 143.615 53.515 144.565 ;
        RECT 53.705 144.530 54.035 145.705 ;
        RECT 54.205 144.905 54.485 145.875 ;
        RECT 53.705 144.380 54.485 144.530 ;
        RECT 55.385 144.380 55.610 146.255 ;
        RECT 55.790 146.245 58.270 146.255 ;
        RECT 58.025 145.480 58.270 146.245 ;
        RECT 57.995 145.170 58.305 145.480 ;
        RECT 58.665 144.995 58.835 147.185 ;
        RECT 60.175 145.925 60.465 147.090 ;
        RECT 61.185 146.285 62.610 146.510 ;
        RECT 60.090 145.755 60.550 145.925 ;
        RECT 59.240 145.375 60.620 145.545 ;
        RECT 59.335 144.995 59.665 145.190 ;
        RECT 58.665 144.825 59.665 144.995 ;
        RECT 53.705 144.155 55.610 144.380 ;
        RECT 59.335 144.405 59.665 144.825 ;
        RECT 59.335 144.235 60.015 144.405 ;
        RECT 60.195 144.235 60.525 145.375 ;
        RECT 53.705 144.000 54.485 144.155 ;
        RECT 59.325 144.050 59.675 144.065 ;
        RECT 53.705 143.495 54.030 144.000 ;
        RECT 59.280 143.855 59.675 144.050 ;
        RECT 54.200 143.325 54.485 143.830 ;
        RECT 59.325 143.815 59.675 143.855 ;
        RECT 59.845 143.635 60.015 144.235 ;
        RECT 60.185 144.055 60.535 144.065 ;
        RECT 61.185 144.055 61.510 146.285 ;
        RECT 65.190 145.375 66.570 145.545 ;
        RECT 65.520 144.575 65.850 145.205 ;
        RECT 63.390 144.210 63.615 144.215 ;
        RECT 65.520 144.210 65.750 144.575 ;
        RECT 66.020 144.555 66.250 145.375 ;
        RECT 60.185 143.830 61.610 144.055 ;
        RECT 63.390 143.995 65.750 144.210 ;
        RECT 63.390 143.990 63.615 143.995 ;
        RECT 65.520 143.975 65.750 143.995 ;
        RECT 60.185 143.815 60.535 143.830 ;
        RECT 53.190 143.155 54.570 143.325 ;
        RECT 59.345 142.825 59.585 143.635 ;
        RECT 59.755 142.995 60.085 143.635 ;
        RECT 60.255 142.825 60.525 143.635 ;
        RECT 65.520 142.995 65.850 143.975 ;
        RECT 66.020 142.825 66.230 143.965 ;
        RECT 66.840 143.275 67.300 143.445 ;
        RECT 59.240 142.655 60.620 142.825 ;
        RECT 65.190 142.655 66.570 142.825 ;
        RECT 66.925 142.110 67.215 143.275 ;
        RECT 49.040 141.175 50.420 141.345 ;
        RECT 49.370 140.375 49.700 141.005 ;
        RECT 49.370 140.365 49.600 140.375 ;
        RECT 48.185 140.135 49.600 140.365 ;
        RECT 49.870 140.355 50.100 141.175 ;
        RECT 66.925 140.725 67.215 141.450 ;
        RECT 66.840 140.555 67.300 140.725 ;
        RECT 49.370 139.775 49.600 140.135 ;
        RECT 49.370 138.795 49.700 139.775 ;
        RECT 49.870 138.625 50.080 139.765 ;
        RECT 50.540 139.025 51.000 139.195 ;
        RECT 49.040 138.455 50.420 138.625 ;
        RECT 50.625 137.860 50.915 139.025 ;
        RECT 44.400 136.525 46.700 136.695 ;
        RECT 44.485 135.805 45.080 136.355 ;
        RECT 45.250 136.125 46.185 136.525 ;
        RECT 50.625 136.475 50.915 137.200 ;
        RECT 68.400 137.135 70.700 137.305 ;
        RECT 68.485 136.565 68.745 136.965 ;
        RECT 68.915 136.735 69.850 137.135 ;
        RECT 70.020 136.625 70.615 136.965 ;
        RECT 70.955 136.665 71.125 136.750 ;
        RECT 73.675 136.665 73.845 136.750 ;
        RECT 46.355 135.955 46.615 136.355 ;
        RECT 50.540 136.305 51.000 136.475 ;
        RECT 68.485 136.395 69.850 136.565 ;
        RECT 44.485 134.655 44.725 135.635 ;
        RECT 44.905 134.485 45.080 135.805 ;
        RECT 45.250 135.785 46.615 135.955 ;
        RECT 45.250 134.715 45.985 135.785 ;
        RECT 46.155 135.540 46.615 135.615 ;
        RECT 46.155 135.355 47.640 135.540 ;
        RECT 46.155 134.885 46.615 135.355 ;
        RECT 47.455 135.295 47.640 135.355 ;
        RECT 69.115 135.325 69.850 136.395 ;
        RECT 48.185 135.295 48.415 135.320 ;
        RECT 47.455 135.110 48.415 135.295 ;
        RECT 48.185 135.090 48.415 135.110 ;
        RECT 68.485 135.155 69.850 135.325 ;
        RECT 70.020 135.305 70.195 136.625 ;
        RECT 70.375 135.810 70.615 136.455 ;
        RECT 70.955 136.375 72.290 136.665 ;
        RECT 72.950 136.375 73.845 136.665 ;
        RECT 70.955 136.290 71.125 136.375 ;
        RECT 73.675 136.290 73.845 136.375 ;
        RECT 70.375 135.770 71.755 135.810 ;
        RECT 70.375 135.595 71.770 135.770 ;
        RECT 70.375 135.475 70.615 135.595 ;
        RECT 68.485 134.755 68.745 135.155 ;
        RECT 45.250 134.545 46.615 134.715 ;
        RECT 68.915 134.585 69.850 134.985 ;
        RECT 70.020 134.755 70.615 135.305 ;
        RECT 44.485 134.145 45.080 134.485 ;
        RECT 45.250 133.975 46.185 134.375 ;
        RECT 46.355 134.145 46.615 134.545 ;
        RECT 46.995 134.375 47.165 134.460 ;
        RECT 49.715 134.375 49.885 134.460 ;
        RECT 68.400 134.415 70.700 134.585 ;
        RECT 46.995 134.085 48.330 134.375 ;
        RECT 48.990 134.085 49.885 134.375 ;
        RECT 46.995 134.000 47.165 134.085 ;
        RECT 49.715 134.000 49.885 134.085 ;
        RECT 44.400 133.805 46.700 133.975 ;
        RECT 71.530 132.130 71.770 135.595 ;
      LAYER mcon ;
        RECT 53.385 161.525 53.555 161.695 ;
        RECT 51.645 159.985 51.815 160.155 ;
        RECT 52.105 159.985 52.275 160.155 ;
        RECT 52.565 159.985 52.735 160.155 ;
        RECT 57.485 159.925 57.655 160.095 ;
        RECT 53.385 158.805 53.555 158.975 ;
        RECT 51.645 157.265 51.815 157.435 ;
        RECT 52.105 157.265 52.275 157.435 ;
        RECT 52.565 157.265 52.735 157.435 ;
        RECT 53.920 157.415 54.090 157.585 ;
        RECT 58.235 158.225 58.405 158.395 ;
        RECT 58.695 158.225 58.865 158.395 ;
        RECT 59.155 158.225 59.325 158.395 ;
        RECT 57.485 157.205 57.655 157.375 ;
        RECT 55.910 156.915 56.095 157.090 ;
        RECT 69.735 157.875 69.905 158.045 ;
        RECT 59.115 157.335 59.285 157.505 ;
        RECT 59.465 156.665 59.635 156.835 ;
        RECT 58.235 155.505 58.405 155.675 ;
        RECT 58.695 155.505 58.865 155.675 ;
        RECT 59.155 155.505 59.325 155.675 ;
        RECT 66.185 155.625 66.355 155.795 ;
        RECT 66.645 155.625 66.815 155.795 ;
        RECT 67.105 155.625 67.275 155.795 ;
        RECT 67.565 155.625 67.735 155.795 ;
        RECT 68.025 155.625 68.195 155.795 ;
        RECT 68.485 155.625 68.655 155.795 ;
        RECT 68.945 155.625 69.115 155.795 ;
        RECT 66.715 154.865 66.885 155.035 ;
        RECT 69.735 155.155 69.905 155.325 ;
        RECT 66.185 152.905 66.355 153.075 ;
        RECT 66.645 152.905 66.815 153.075 ;
        RECT 67.105 152.905 67.275 153.075 ;
        RECT 67.565 152.905 67.735 153.075 ;
        RECT 68.025 152.905 68.195 153.075 ;
        RECT 68.485 152.905 68.655 153.075 ;
        RECT 68.945 152.905 69.115 153.075 ;
        RECT 59.465 151.515 59.635 151.685 ;
        RECT 59.465 151.055 59.635 151.225 ;
        RECT 61.365 151.325 61.635 151.595 ;
        RECT 62.185 151.515 62.355 151.685 ;
        RECT 62.185 151.055 62.355 151.225 ;
        RECT 61.010 150.810 61.190 150.990 ;
        RECT 59.465 150.595 59.635 150.765 ;
        RECT 62.185 150.595 62.355 150.765 ;
        RECT 57.405 149.835 57.575 150.005 ;
        RECT 60.125 149.835 60.295 150.005 ;
        RECT 60.235 148.475 60.405 148.645 ;
        RECT 52.685 147.425 52.855 147.595 ;
        RECT 58.665 147.015 58.835 147.185 ;
        RECT 53.335 145.875 53.505 146.045 ;
        RECT 53.795 145.875 53.965 146.045 ;
        RECT 54.255 145.875 54.425 146.045 ;
        RECT 52.685 144.705 52.855 144.875 ;
        RECT 62.415 146.315 62.585 146.485 ;
        RECT 60.235 145.755 60.405 145.925 ;
        RECT 59.385 145.375 59.555 145.545 ;
        RECT 59.845 145.375 60.015 145.545 ;
        RECT 60.305 145.375 60.475 145.545 ;
        RECT 59.280 143.855 59.475 144.050 ;
        RECT 65.335 145.375 65.505 145.545 ;
        RECT 65.795 145.375 65.965 145.545 ;
        RECT 66.255 145.375 66.425 145.545 ;
        RECT 53.335 143.155 53.505 143.325 ;
        RECT 53.795 143.155 53.965 143.325 ;
        RECT 54.255 143.155 54.425 143.325 ;
        RECT 66.985 143.275 67.155 143.445 ;
        RECT 59.385 142.655 59.555 142.825 ;
        RECT 59.845 142.655 60.015 142.825 ;
        RECT 60.305 142.655 60.475 142.825 ;
        RECT 65.335 142.655 65.505 142.825 ;
        RECT 65.795 142.655 65.965 142.825 ;
        RECT 66.255 142.655 66.425 142.825 ;
        RECT 49.185 141.175 49.355 141.345 ;
        RECT 49.645 141.175 49.815 141.345 ;
        RECT 50.105 141.175 50.275 141.345 ;
        RECT 66.985 140.555 67.155 140.725 ;
        RECT 50.685 139.025 50.855 139.195 ;
        RECT 49.185 138.455 49.355 138.625 ;
        RECT 49.645 138.455 49.815 138.625 ;
        RECT 50.105 138.455 50.275 138.625 ;
        RECT 44.545 136.525 44.715 136.695 ;
        RECT 45.005 136.525 45.175 136.695 ;
        RECT 45.465 136.525 45.635 136.695 ;
        RECT 45.925 136.525 46.095 136.695 ;
        RECT 46.385 136.525 46.555 136.695 ;
        RECT 44.485 135.975 44.655 136.145 ;
        RECT 68.545 137.135 68.715 137.305 ;
        RECT 69.005 137.135 69.175 137.305 ;
        RECT 69.465 137.135 69.635 137.305 ;
        RECT 69.925 137.135 70.095 137.305 ;
        RECT 70.385 137.135 70.555 137.305 ;
        RECT 50.685 136.305 50.855 136.475 ;
        RECT 44.485 135.125 44.725 135.365 ;
        RECT 70.955 136.435 71.125 136.605 ;
        RECT 73.675 136.435 73.845 136.605 ;
        RECT 68.545 134.415 68.715 134.585 ;
        RECT 69.005 134.415 69.175 134.585 ;
        RECT 69.465 134.415 69.635 134.585 ;
        RECT 69.925 134.415 70.095 134.585 ;
        RECT 70.385 134.415 70.555 134.585 ;
        RECT 46.995 134.145 47.165 134.315 ;
        RECT 49.715 134.145 49.885 134.315 ;
        RECT 44.545 133.805 44.715 133.975 ;
        RECT 45.005 133.805 45.175 133.975 ;
        RECT 45.465 133.805 45.635 133.975 ;
        RECT 45.925 133.805 46.095 133.975 ;
        RECT 46.385 133.805 46.555 133.975 ;
      LAYER met1 ;
        RECT 50.125 162.420 53.625 162.575 ;
        RECT 50.125 153.825 50.280 162.420 ;
        RECT 53.470 161.850 53.625 162.420 ;
        RECT 53.240 161.825 55.625 161.850 ;
        RECT 52.625 161.815 55.625 161.825 ;
        RECT 52.575 161.695 55.625 161.815 ;
        RECT 52.575 161.670 53.700 161.695 ;
        RECT 52.575 161.495 52.835 161.670 ;
        RECT 53.240 161.370 53.700 161.670 ;
        RECT 55.470 160.380 55.625 161.695 ;
        RECT 50.725 160.310 51.575 160.325 ;
        RECT 50.725 160.300 52.880 160.310 ;
        RECT 50.725 160.170 53.170 160.300 ;
        RECT 55.470 160.225 68.725 160.380 ;
        RECT 50.725 154.775 50.880 160.170 ;
        RECT 51.500 160.160 53.170 160.170 ;
        RECT 51.500 159.830 52.880 160.160 ;
        RECT 53.030 159.570 53.170 160.160 ;
        RECT 57.340 159.770 57.800 160.225 ;
        RECT 52.880 159.430 53.170 159.570 ;
        RECT 61.070 159.670 65.775 159.825 ;
        RECT 52.880 159.120 53.020 159.430 ;
        RECT 53.240 159.120 53.700 159.130 ;
        RECT 52.880 158.980 53.700 159.120 ;
        RECT 53.240 158.795 53.700 158.980 ;
        RECT 53.240 158.655 55.320 158.795 ;
        RECT 61.070 158.775 61.225 159.670 ;
        RECT 53.240 158.650 53.700 158.655 ;
        RECT 51.500 157.110 52.880 157.590 ;
        RECT 53.890 157.355 54.120 157.645 ;
        RECT 55.180 157.470 55.320 158.655 ;
        RECT 59.315 158.620 61.225 158.775 ;
        RECT 61.790 159.130 65.295 159.420 ;
        RECT 59.315 158.550 59.470 158.620 ;
        RECT 57.725 158.395 59.470 158.550 ;
        RECT 57.725 157.930 57.880 158.395 ;
        RECT 58.090 158.070 59.470 158.395 ;
        RECT 57.725 157.775 58.075 157.930 ;
        RECT 57.920 157.620 58.075 157.775 ;
        RECT 57.735 157.530 58.115 157.620 ;
        RECT 51.525 156.965 51.680 157.110 ;
        RECT 51.475 156.645 51.735 156.965 ;
        RECT 52.680 155.680 52.835 157.110 ;
        RECT 53.915 157.090 54.090 157.355 ;
        RECT 55.180 157.330 56.620 157.470 ;
        RECT 56.480 157.170 56.620 157.330 ;
        RECT 57.340 157.385 58.115 157.530 ;
        RECT 59.085 157.505 59.315 157.535 ;
        RECT 61.790 157.505 62.080 159.130 ;
        RECT 57.340 157.170 57.800 157.385 ;
        RECT 59.045 157.335 62.085 157.505 ;
        RECT 59.085 157.305 59.315 157.335 ;
        RECT 55.850 157.090 56.155 157.120 ;
        RECT 53.910 156.915 56.155 157.090 ;
        RECT 56.480 157.050 57.800 157.170 ;
        RECT 56.480 157.030 57.420 157.050 ;
        RECT 55.850 156.885 56.155 156.915 ;
        RECT 59.405 156.840 59.695 156.865 ;
        RECT 59.405 156.805 61.040 156.840 ;
        RECT 59.405 156.660 61.055 156.805 ;
        RECT 59.405 156.635 59.695 156.660 ;
        RECT 52.680 155.525 57.675 155.680 ;
        RECT 57.520 155.380 57.675 155.525 ;
        RECT 58.090 155.475 59.470 155.830 ;
        RECT 58.020 155.385 59.470 155.475 ;
        RECT 58.020 155.380 60.375 155.385 ;
        RECT 57.520 155.230 60.375 155.380 ;
        RECT 57.520 155.225 58.175 155.230 ;
        RECT 50.725 154.620 59.465 154.775 ;
        RECT 50.125 153.670 57.405 153.825 ;
        RECT 57.250 150.150 57.405 153.670 ;
        RECT 59.310 151.830 59.465 154.620 ;
        RECT 60.220 152.885 60.375 155.230 ;
        RECT 60.845 153.605 61.055 156.660 ;
        RECT 65.005 154.235 65.295 159.130 ;
        RECT 65.620 156.230 65.775 159.670 ;
        RECT 68.570 158.230 68.725 160.225 ;
        RECT 68.570 158.075 75.075 158.230 ;
        RECT 69.590 157.720 70.050 158.075 ;
        RECT 65.620 156.075 66.425 156.230 ;
        RECT 65.975 155.950 66.425 156.075 ;
        RECT 65.975 155.925 69.260 155.950 ;
        RECT 66.040 155.675 69.260 155.925 ;
        RECT 66.040 155.575 69.330 155.675 ;
        RECT 66.040 155.470 69.430 155.575 ;
        RECT 69.175 155.420 69.430 155.470 ;
        RECT 69.275 155.155 69.430 155.420 ;
        RECT 69.590 155.155 70.050 155.480 ;
        RECT 65.540 155.035 65.860 155.130 ;
        RECT 69.275 155.080 70.050 155.155 ;
        RECT 70.375 155.080 73.525 155.175 ;
        RECT 66.655 155.035 66.945 155.065 ;
        RECT 65.540 154.870 66.945 155.035 ;
        RECT 69.275 155.020 73.525 155.080 ;
        RECT 69.275 155.000 70.530 155.020 ;
        RECT 69.925 154.925 70.530 155.000 ;
        RECT 65.615 154.865 66.945 154.870 ;
        RECT 66.655 154.835 66.945 154.865 ;
        RECT 66.850 154.235 67.080 154.295 ;
        RECT 65.005 154.065 67.080 154.235 ;
        RECT 65.005 154.055 65.295 154.065 ;
        RECT 66.850 154.005 67.080 154.065 ;
        RECT 60.845 153.585 62.655 153.605 ;
        RECT 60.845 153.395 62.665 153.585 ;
        RECT 70.095 153.525 70.415 153.785 ;
        RECT 62.335 153.325 62.665 153.395 ;
        RECT 66.040 152.925 69.260 153.230 ;
        RECT 70.125 152.925 70.280 153.525 ;
        RECT 60.220 152.730 62.675 152.885 ;
        RECT 61.365 152.515 61.985 152.535 ;
        RECT 61.365 152.265 62.085 152.515 ;
        RECT 59.310 150.450 59.790 151.830 ;
        RECT 61.365 151.655 61.635 152.265 ;
        RECT 61.815 152.185 62.085 152.265 ;
        RECT 62.520 151.930 62.675 152.730 ;
        RECT 62.325 151.830 62.675 151.930 ;
        RECT 62.030 151.775 62.675 151.830 ;
        RECT 64.670 152.770 70.575 152.925 ;
        RECT 61.335 151.265 61.665 151.655 ;
        RECT 61.010 151.020 61.190 151.090 ;
        RECT 60.950 150.780 61.250 151.020 ;
        RECT 61.010 150.620 61.190 150.780 ;
        RECT 60.930 150.560 61.190 150.620 ;
        RECT 62.030 150.605 62.510 151.775 ;
        RECT 64.670 150.605 64.825 152.770 ;
        RECT 66.040 152.750 69.260 152.770 ;
        RECT 65.570 152.240 65.830 152.560 ;
        RECT 65.615 151.335 65.785 152.240 ;
        RECT 65.615 151.165 70.215 151.335 ;
        RECT 59.310 150.230 59.465 150.450 ;
        RECT 59.310 150.150 60.125 150.230 ;
        RECT 55.745 150.025 56.065 150.080 ;
        RECT 57.250 150.025 57.730 150.150 ;
        RECT 59.310 150.075 60.450 150.150 ;
        RECT 55.745 149.870 57.730 150.025 ;
        RECT 55.745 149.820 56.065 149.870 ;
        RECT 57.250 149.690 57.730 149.870 ;
        RECT 59.970 149.690 60.450 150.075 ;
        RECT 47.525 149.530 50.180 149.675 ;
        RECT 60.295 149.530 60.450 149.690 ;
        RECT 47.525 149.520 60.450 149.530 ;
        RECT 47.525 146.780 47.680 149.520 ;
        RECT 50.025 149.375 60.450 149.520 ;
        RECT 49.440 149.220 49.760 149.230 ;
        RECT 60.930 149.220 61.170 150.560 ;
        RECT 49.440 148.980 61.170 149.220 ;
        RECT 62.030 150.450 64.825 150.605 ;
        RECT 49.440 148.970 49.760 148.980 ;
        RECT 53.025 148.780 60.550 148.800 ;
        RECT 62.030 148.780 62.185 150.450 ;
        RECT 53.025 148.645 62.185 148.780 ;
        RECT 53.025 147.930 53.180 148.645 ;
        RECT 60.090 148.625 62.185 148.645 ;
        RECT 60.090 148.320 60.550 148.625 ;
        RECT 55.775 147.930 56.035 148.110 ;
        RECT 50.195 147.825 50.515 147.880 ;
        RECT 53.025 147.830 56.035 147.930 ;
        RECT 50.195 147.750 52.675 147.825 ;
        RECT 52.875 147.790 56.035 147.830 ;
        RECT 52.875 147.775 55.980 147.790 ;
        RECT 52.875 147.750 53.180 147.775 ;
        RECT 50.195 147.675 53.180 147.750 ;
        RECT 50.195 147.670 53.000 147.675 ;
        RECT 50.195 147.620 50.515 147.670 ;
        RECT 52.540 147.270 53.000 147.670 ;
        RECT 58.605 147.185 58.895 147.215 ;
        RECT 70.045 147.185 70.215 151.165 ;
        RECT 58.605 147.015 70.215 147.185 ;
        RECT 58.605 146.985 58.895 147.015 ;
        RECT 47.525 146.625 51.320 146.780 ;
        RECT 51.130 144.680 51.285 146.625 ;
        RECT 54.525 146.620 58.680 146.775 ;
        RECT 54.525 146.280 54.680 146.620 ;
        RECT 54.425 146.200 54.680 146.280 ;
        RECT 53.190 146.125 54.680 146.200 ;
        RECT 58.525 146.125 58.680 146.620 ;
        RECT 62.355 146.510 62.645 146.515 ;
        RECT 62.355 146.285 63.610 146.510 ;
        RECT 69.540 146.425 69.860 146.480 ;
        RECT 53.190 145.875 54.570 146.125 ;
        RECT 58.525 145.970 59.425 146.125 ;
        RECT 53.020 145.720 54.570 145.875 ;
        RECT 53.020 145.030 53.175 145.720 ;
        RECT 59.270 145.700 59.425 145.970 ;
        RECT 60.090 145.700 60.550 146.080 ;
        RECT 59.240 145.545 62.225 145.700 ;
        RECT 57.935 145.140 58.365 145.510 ;
        RECT 59.240 145.220 60.620 145.545 ;
        RECT 52.540 144.875 53.175 145.030 ;
        RECT 52.540 144.680 53.000 144.875 ;
        RECT 51.130 144.550 53.000 144.680 ;
        RECT 51.130 144.525 52.875 144.550 ;
        RECT 49.440 144.120 49.760 144.130 ;
        RECT 39.150 143.880 53.515 144.120 ;
        RECT 57.995 144.050 58.305 145.140 ;
        RECT 59.250 144.050 59.505 144.080 ;
        RECT 39.150 138.420 39.390 143.880 ;
        RECT 49.440 143.870 49.760 143.880 ;
        RECT 57.995 143.855 59.545 144.050 ;
        RECT 57.995 143.845 58.305 143.855 ;
        RECT 59.250 143.825 59.505 143.855 ;
        RECT 50.175 143.155 50.435 143.240 ;
        RECT 53.190 143.155 54.570 143.480 ;
        RECT 50.175 143.000 54.570 143.155 ;
        RECT 50.175 142.920 50.435 143.000 ;
        RECT 51.570 141.500 51.725 143.000 ;
        RECT 54.375 142.655 54.530 143.000 ;
        RECT 59.240 142.655 60.620 142.980 ;
        RECT 54.375 142.500 60.620 142.655 ;
        RECT 62.070 142.860 62.225 145.545 ;
        RECT 63.385 144.275 63.610 146.285 ;
        RECT 64.320 146.270 69.860 146.425 ;
        RECT 63.360 143.930 63.645 144.275 ;
        RECT 63.385 143.890 63.610 143.930 ;
        RECT 64.320 143.030 64.475 146.270 ;
        RECT 69.540 146.220 69.860 146.270 ;
        RECT 66.375 145.700 67.080 145.775 ;
        RECT 64.825 145.620 67.080 145.700 ;
        RECT 64.825 145.545 66.570 145.620 ;
        RECT 62.070 142.540 62.330 142.860 ;
        RECT 64.240 142.770 64.560 143.030 ;
        RECT 64.320 142.630 64.475 142.770 ;
        RECT 60.275 142.080 60.430 142.500 ;
        RECT 64.825 142.080 64.980 145.545 ;
        RECT 65.190 145.220 66.570 145.545 ;
        RECT 66.925 145.530 67.080 145.620 ;
        RECT 70.420 145.530 70.575 152.770 ;
        RECT 72.295 146.425 72.615 146.480 ;
        RECT 73.370 146.425 73.525 155.020 ;
        RECT 74.920 153.815 75.075 158.075 ;
        RECT 74.870 153.495 75.130 153.815 ;
        RECT 72.295 146.270 73.525 146.425 ;
        RECT 72.295 146.220 72.615 146.270 ;
        RECT 66.925 145.375 70.575 145.530 ;
        RECT 67.125 143.600 68.480 143.675 ;
        RECT 66.840 143.520 68.480 143.600 ;
        RECT 66.840 143.275 67.300 143.520 ;
        RECT 66.770 143.120 67.300 143.275 ;
        RECT 65.190 142.655 66.570 142.980 ;
        RECT 66.770 142.655 66.925 143.120 ;
        RECT 65.190 142.500 66.925 142.655 ;
        RECT 60.275 141.925 64.980 142.080 ;
        RECT 46.575 141.345 51.725 141.500 ;
        RECT 39.150 138.180 43.720 138.420 ;
        RECT 43.515 136.145 43.685 138.180 ;
        RECT 46.575 136.850 46.730 141.345 ;
        RECT 49.040 141.020 50.420 141.345 ;
        RECT 64.245 141.080 64.565 141.135 ;
        RECT 65.670 141.080 65.825 142.500 ;
        RECT 64.245 140.925 65.825 141.080 ;
        RECT 64.245 140.875 64.565 140.925 ;
        RECT 44.175 136.775 46.730 136.850 ;
        RECT 47.575 140.720 48.875 140.875 ;
        RECT 62.040 140.770 62.360 140.825 ;
        RECT 44.175 136.695 46.700 136.775 ;
        RECT 44.400 136.370 46.700 136.695 ;
        RECT 44.455 136.145 44.685 136.175 ;
        RECT 43.515 135.975 45.080 136.145 ;
        RECT 44.455 135.945 44.685 135.975 ;
        RECT 43.480 135.365 43.720 135.370 ;
        RECT 44.455 135.365 44.755 135.425 ;
        RECT 43.480 135.125 44.755 135.365 ;
        RECT 43.480 132.370 43.720 135.125 ;
        RECT 44.455 135.065 44.755 135.125 ;
        RECT 47.575 134.930 47.730 140.720 ;
        RECT 48.155 140.075 48.445 140.425 ;
        RECT 48.185 135.380 48.415 140.075 ;
        RECT 48.720 138.430 48.875 140.720 ;
        RECT 50.675 140.615 62.360 140.770 ;
        RECT 50.675 139.775 50.830 140.615 ;
        RECT 62.040 140.565 62.360 140.615 ;
        RECT 66.840 140.555 67.300 140.880 ;
        RECT 63.425 140.400 67.300 140.555 ;
        RECT 50.675 139.620 51.000 139.775 ;
        RECT 50.845 139.350 51.000 139.620 ;
        RECT 50.540 139.025 51.000 139.350 ;
        RECT 63.425 139.280 63.580 140.400 ;
        RECT 50.375 138.870 51.000 139.025 ;
        RECT 63.345 139.020 63.665 139.280 ;
        RECT 67.130 139.180 67.285 140.400 ;
        RECT 68.325 140.025 68.480 143.520 ;
        RECT 70.090 140.025 70.410 140.080 ;
        RECT 68.325 139.870 70.410 140.025 ;
        RECT 70.090 139.820 70.410 139.870 ;
        RECT 71.720 139.790 71.980 140.110 ;
        RECT 67.125 139.160 67.285 139.180 ;
        RECT 63.425 138.975 63.580 139.020 ;
        RECT 50.375 138.830 50.530 138.870 ;
        RECT 67.075 138.840 67.335 139.160 ;
        RECT 50.275 138.780 50.530 138.830 ;
        RECT 49.040 138.675 50.530 138.780 ;
        RECT 49.040 138.430 50.420 138.675 ;
        RECT 48.720 138.300 50.420 138.430 ;
        RECT 48.720 138.275 50.325 138.300 ;
        RECT 71.770 137.460 71.925 139.790 ;
        RECT 73.570 138.890 73.830 139.210 ;
        RECT 68.400 137.305 71.925 137.460 ;
        RECT 73.620 137.430 73.775 138.890 ;
        RECT 68.400 137.125 70.700 137.305 ;
        RECT 73.620 137.275 74.025 137.430 ;
        RECT 68.400 136.980 70.955 137.125 ;
        RECT 70.575 136.970 70.955 136.980 ;
        RECT 70.800 136.750 70.955 136.970 ;
        RECT 73.870 136.750 74.025 137.275 ;
        RECT 50.540 136.275 51.000 136.630 ;
        RECT 70.800 136.425 71.280 136.750 ;
        RECT 49.885 136.150 51.000 136.275 ;
        RECT 49.885 136.120 50.675 136.150 ;
        RECT 48.155 135.030 48.445 135.380 ;
        RECT 46.825 134.775 47.730 134.930 ;
        RECT 46.825 134.460 46.980 134.775 ;
        RECT 49.885 134.460 50.040 136.120 ;
        RECT 50.845 135.030 51.000 136.150 ;
        RECT 70.775 136.290 71.280 136.425 ;
        RECT 73.520 136.675 74.025 136.750 ;
        RECT 73.520 136.425 74.000 136.675 ;
        RECT 73.520 136.290 74.225 136.425 ;
        RECT 70.775 135.975 70.930 136.290 ;
        RECT 73.875 136.270 74.225 136.290 ;
        RECT 70.775 135.820 71.025 135.975 ;
        RECT 74.070 135.825 74.225 136.270 ;
        RECT 63.345 135.030 63.665 135.085 ;
        RECT 50.845 134.875 66.225 135.030 ;
        RECT 63.345 134.825 63.665 134.875 ;
        RECT 46.825 134.180 47.320 134.460 ;
        RECT 46.525 134.130 47.320 134.180 ;
        RECT 44.400 134.025 47.320 134.130 ;
        RECT 44.400 133.725 46.700 134.025 ;
        RECT 46.840 134.000 47.320 134.025 ;
        RECT 49.560 134.235 50.040 134.460 ;
        RECT 66.070 134.380 66.225 134.875 ;
        RECT 68.400 134.380 70.700 134.740 ;
        RECT 51.070 134.235 51.330 134.315 ;
        RECT 49.560 134.080 51.330 134.235 ;
        RECT 66.070 134.260 70.700 134.380 ;
        RECT 66.070 134.225 68.675 134.260 ;
        RECT 49.560 134.000 50.040 134.080 ;
        RECT 51.070 133.995 51.330 134.080 ;
        RECT 69.845 134.020 70.165 134.260 ;
        RECT 69.925 133.975 70.080 134.020 ;
        RECT 47.525 133.725 47.785 133.810 ;
        RECT 70.870 133.725 71.025 135.820 ;
        RECT 44.400 133.650 71.025 133.725 ;
        RECT 46.430 133.570 71.025 133.650 ;
        RECT 73.070 135.670 74.225 135.825 ;
        RECT 47.525 133.490 47.785 133.570 ;
        RECT 71.470 132.370 71.830 132.400 ;
        RECT 43.480 132.130 71.830 132.370 ;
        RECT 71.470 132.100 71.830 132.130 ;
        RECT 73.070 132.115 73.225 135.670 ;
        RECT 47.525 131.640 47.785 131.960 ;
        RECT 73.020 131.795 73.280 132.115 ;
        RECT 47.575 129.680 47.730 131.640 ;
        RECT 2.425 129.525 47.730 129.680 ;
      LAYER via ;
        RECT 52.575 161.525 52.835 161.785 ;
        RECT 51.475 156.675 51.735 156.935 ;
        RECT 65.570 154.870 65.830 155.130 ;
        RECT 62.365 153.325 62.635 153.585 ;
        RECT 70.125 153.525 70.385 153.785 ;
        RECT 61.815 152.215 62.085 152.485 ;
        RECT 65.570 152.270 65.830 152.530 ;
        RECT 55.775 149.820 56.035 150.080 ;
        RECT 49.470 148.970 49.730 149.230 ;
        RECT 50.225 147.620 50.485 147.880 ;
        RECT 55.775 147.820 56.035 148.080 ;
        RECT 49.470 143.870 49.730 144.130 ;
        RECT 50.175 142.950 50.435 143.210 ;
        RECT 69.570 146.220 69.830 146.480 ;
        RECT 62.070 142.570 62.330 142.830 ;
        RECT 64.270 142.770 64.530 143.030 ;
        RECT 72.325 146.220 72.585 146.480 ;
        RECT 74.870 153.525 75.130 153.785 ;
        RECT 64.275 140.875 64.535 141.135 ;
        RECT 62.070 140.565 62.330 140.825 ;
        RECT 63.375 139.020 63.635 139.280 ;
        RECT 70.120 139.820 70.380 140.080 ;
        RECT 71.720 139.820 71.980 140.080 ;
        RECT 67.075 138.870 67.335 139.130 ;
        RECT 73.570 138.920 73.830 139.180 ;
        RECT 63.375 134.825 63.635 135.085 ;
        RECT 51.070 134.025 51.330 134.285 ;
        RECT 69.875 134.020 70.135 134.280 ;
        RECT 47.525 133.520 47.785 133.780 ;
        RECT 47.525 131.670 47.785 131.930 ;
        RECT 73.020 131.825 73.280 132.085 ;
      LAYER met2 ;
        RECT 52.625 161.785 52.780 161.825 ;
        RECT 52.545 161.525 52.865 161.785 ;
        RECT 52.625 160.575 52.780 161.525 ;
        RECT 52.625 160.420 54.825 160.575 ;
        RECT 51.445 156.675 51.765 156.935 ;
        RECT 51.525 155.880 51.680 156.675 ;
        RECT 54.670 155.880 54.825 160.420 ;
        RECT 51.525 155.725 54.825 155.880 ;
        RECT 65.570 154.840 65.830 155.160 ;
        RECT 62.365 152.485 62.635 153.615 ;
        RECT 65.615 152.530 65.785 154.840 ;
        RECT 70.125 153.730 70.385 153.815 ;
        RECT 74.840 153.730 75.160 153.785 ;
        RECT 70.125 153.575 75.160 153.730 ;
        RECT 70.125 153.495 70.385 153.575 ;
        RECT 74.840 153.525 75.160 153.575 ;
        RECT 61.785 152.215 62.635 152.485 ;
        RECT 65.540 152.270 65.860 152.530 ;
        RECT 55.775 149.790 56.035 150.110 ;
        RECT 49.470 148.940 49.730 149.260 ;
        RECT 49.480 144.160 49.720 148.940 ;
        RECT 55.825 148.080 55.980 149.790 ;
        RECT 50.225 147.590 50.485 147.910 ;
        RECT 55.745 147.820 56.065 148.080 ;
        RECT 55.825 147.775 55.980 147.820 ;
        RECT 49.470 143.840 49.730 144.160 ;
        RECT 50.225 143.210 50.380 147.590 ;
        RECT 69.570 146.425 69.830 146.510 ;
        RECT 72.325 146.425 72.585 146.510 ;
        RECT 69.570 146.270 72.585 146.425 ;
        RECT 69.570 146.190 69.830 146.270 ;
        RECT 72.325 146.190 72.585 146.270 ;
        RECT 50.145 142.950 50.465 143.210 ;
        RECT 62.040 142.570 62.360 142.830 ;
        RECT 64.270 142.740 64.530 143.060 ;
        RECT 62.120 140.855 62.275 142.570 ;
        RECT 64.320 141.165 64.475 142.740 ;
        RECT 62.070 140.535 62.330 140.855 ;
        RECT 64.275 140.845 64.535 141.165 ;
        RECT 70.120 140.025 70.380 140.110 ;
        RECT 71.690 140.025 72.010 140.080 ;
        RECT 70.120 139.870 72.010 140.025 ;
        RECT 70.120 139.790 70.380 139.870 ;
        RECT 71.690 139.820 72.010 139.870 ;
        RECT 63.375 138.990 63.635 139.310 ;
        RECT 67.045 139.080 67.365 139.130 ;
        RECT 73.540 139.080 73.860 139.180 ;
        RECT 42.325 136.695 44.330 136.850 ;
        RECT 42.325 134.335 42.480 136.695 ;
        RECT 63.425 135.115 63.580 138.990 ;
        RECT 67.045 138.925 73.860 139.080 ;
        RECT 67.045 138.870 67.365 138.925 ;
        RECT 73.540 138.920 73.860 138.925 ;
        RECT 63.375 134.795 63.635 135.115 ;
        RECT 10.575 134.180 42.480 134.335 ;
        RECT 42.325 131.230 42.480 134.180 ;
        RECT 51.040 134.025 51.360 134.285 ;
        RECT 47.495 133.520 47.815 133.780 ;
        RECT 47.575 131.930 47.730 133.520 ;
        RECT 47.495 131.670 47.815 131.930 ;
        RECT 47.575 131.625 47.730 131.670 ;
        RECT 51.120 131.230 51.275 134.025 ;
        RECT 69.875 133.990 70.135 134.310 ;
        RECT 69.925 132.030 70.080 133.990 ;
        RECT 72.990 132.030 73.310 132.085 ;
        RECT 69.925 131.875 73.310 132.030 ;
        RECT 71.820 131.230 71.975 131.875 ;
        RECT 72.990 131.825 73.310 131.875 ;
        RECT 42.325 131.075 71.975 131.230 ;
        RECT 2.425 129.525 2.580 130.225 ;
  END
END tt_um_test_5
END LIBRARY

