VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_template
  CLASS BLOCK ;
  FOREIGN tt_um_template ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 54.560 209.800 55.155 209.805 ;
        RECT 54.560 209.465 56.165 209.800 ;
        RECT 54.560 208.145 54.735 209.465 ;
        RECT 54.560 207.595 55.155 208.145 ;
      LAYER mcon ;
        RECT 55.910 209.545 56.080 209.715 ;
      LAYER met1 ;
        RECT 55.830 215.930 66.715 216.075 ;
        RECT 55.830 215.740 66.725 215.930 ;
        RECT 55.830 209.830 56.165 215.740 ;
        RECT 66.365 214.920 66.725 215.740 ;
        RECT 55.800 209.435 56.195 209.830 ;
        RECT 55.830 209.385 56.165 209.435 ;
      LAYER via ;
        RECT 66.415 215.020 66.675 215.280 ;
      LAYER met2 ;
        RECT 66.360 23.315 66.735 215.435 ;
        RECT 150.345 23.315 152.475 23.380 ;
        RECT 66.360 22.940 152.475 23.315 ;
        RECT 150.345 22.870 152.475 22.940 ;
      LAYER via2 ;
        RECT 151.950 22.940 152.325 23.315 ;
      LAYER met3 ;
        RECT 151.690 0.280 152.590 23.445 ;
      LAYER via3 ;
        RECT 151.960 0.380 152.400 0.860 ;
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 25.190 197.255 26.390 197.495 ;
      LAYER mcon ;
        RECT 25.280 197.310 25.450 197.480 ;
      LAYER met1 ;
        RECT 21.305 200.755 25.490 201.005 ;
        RECT 20.540 199.475 20.860 199.480 ;
        RECT 21.305 199.475 21.555 200.755 ;
        RECT 20.540 199.225 21.555 199.475 ;
        RECT 20.540 199.220 20.860 199.225 ;
        RECT 25.240 197.245 25.490 200.755 ;
      LAYER via ;
        RECT 20.570 199.220 20.830 199.480 ;
      LAYER met2 ;
        RECT 20.570 199.190 20.830 199.510 ;
        RECT 20.575 26.875 20.825 199.190 ;
        RECT 35.625 26.875 36.575 26.880 ;
        RECT 20.575 26.625 36.575 26.875 ;
        RECT 35.960 25.760 36.545 26.625 ;
      LAYER via2 ;
        RECT 36.110 25.910 36.390 26.190 ;
      LAYER met3 ;
        RECT 35.970 13.470 36.530 26.330 ;
        RECT 35.970 12.910 133.340 13.470 ;
        RECT 132.780 0.130 133.340 12.910 ;
      LAYER via3 ;
        RECT 132.890 0.160 133.240 0.570 ;
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 24.850 213.395 25.315 213.445 ;
        RECT 24.850 213.185 25.950 213.395 ;
        RECT 24.850 213.140 25.315 213.185 ;
        RECT 25.620 213.155 25.950 213.185 ;
      LAYER mcon ;
        RECT 24.905 213.235 25.075 213.405 ;
      LAYER met1 ;
        RECT 10.985 216.905 11.765 216.945 ;
        RECT 10.985 216.655 24.455 216.905 ;
        RECT 10.985 216.615 11.765 216.655 ;
        RECT 24.205 213.445 24.455 216.655 ;
        RECT 24.840 213.445 25.145 213.475 ;
        RECT 24.205 213.195 25.345 213.445 ;
        RECT 24.840 213.170 25.145 213.195 ;
      LAYER via ;
        RECT 11.120 216.650 11.380 216.910 ;
      LAYER met2 ;
        RECT 11.095 13.260 11.410 216.955 ;
        RECT 11.095 12.945 17.205 13.260 ;
        RECT 16.890 7.730 17.205 12.945 ;
        RECT 16.865 6.920 17.225 7.730 ;
      LAYER via2 ;
        RECT 16.905 7.015 17.185 7.295 ;
      LAYER met3 ;
        RECT 16.800 7.400 113.955 7.410 ;
        RECT 16.800 6.920 114.120 7.400 ;
        RECT 113.115 0.180 114.120 6.920 ;
      LAYER via3 ;
        RECT 113.350 0.510 113.840 0.890 ;
      LAYER met4 ;
        RECT 113.170 0.985 114.065 0.995 ;
        RECT 113.170 0.000 114.070 0.985 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 0.223500 ;
    ANTENNADIFFAREA 5.549500 ;
    PORT
      LAYER nwell ;
        RECT 30.910 216.000 33.750 216.010 ;
        RECT 23.250 214.990 24.090 215.000 ;
        RECT 23.250 213.395 26.870 214.990 ;
        RECT 30.910 214.405 34.125 216.000 ;
        RECT 33.285 214.395 34.125 214.405 ;
        RECT 23.900 213.385 26.870 213.395 ;
        RECT 23.900 209.095 27.010 210.700 ;
        RECT 41.150 208.695 46.340 210.300 ;
        RECT 52.750 208.645 57.140 210.250 ;
        RECT 33.900 205.380 34.740 205.400 ;
        RECT 24.270 205.330 27.130 205.350 ;
        RECT 23.960 203.745 27.130 205.330 ;
        RECT 31.260 203.795 34.740 205.380 ;
        RECT 31.260 203.775 34.200 203.795 ;
        RECT 23.960 203.725 24.800 203.745 ;
        RECT 55.460 199.600 58.200 199.610 ;
        RECT 24.290 197.485 27.310 199.090 ;
        RECT 55.460 198.005 58.840 199.600 ;
        RECT 58.000 197.995 58.840 198.005 ;
        RECT 49.530 192.100 50.370 192.120 ;
        RECT 46.300 190.515 50.370 192.100 ;
        RECT 46.300 190.495 50.030 190.515 ;
      LAYER li1 ;
        RECT 31.100 215.735 32.480 215.905 ;
        RECT 23.440 214.725 23.900 214.895 ;
        RECT 23.525 213.560 23.815 214.725 ;
        RECT 25.300 214.715 26.680 214.885 ;
        RECT 25.640 213.575 25.850 214.715 ;
        RECT 32.055 214.595 32.385 215.735 ;
        RECT 33.475 215.725 33.935 215.895 ;
        RECT 33.560 214.560 33.850 215.725 ;
        RECT 24.090 210.425 24.550 210.595 ;
        RECT 25.440 210.425 26.820 210.595 ;
        RECT 24.175 209.260 24.465 210.425 ;
        RECT 25.780 209.285 25.990 210.425 ;
        RECT 41.340 210.025 44.560 210.195 ;
        RECT 45.690 210.025 46.150 210.195 ;
        RECT 42.395 209.175 42.565 210.025 ;
        RECT 43.235 209.515 43.405 210.025 ;
        RECT 45.775 208.860 46.065 210.025 ;
        RECT 52.940 209.975 55.240 210.145 ;
        RECT 56.490 209.975 56.950 210.145 ;
        RECT 53.455 209.575 54.390 209.975 ;
        RECT 56.575 208.810 56.865 209.975 ;
        RECT 24.150 205.055 24.610 205.225 ;
        RECT 25.560 205.075 26.940 205.245 ;
        RECT 31.450 205.105 32.830 205.275 ;
        RECT 34.090 205.125 34.550 205.295 ;
        RECT 24.235 203.890 24.525 205.055 ;
        RECT 25.900 203.935 26.110 205.075 ;
        RECT 32.405 203.965 32.735 205.105 ;
        RECT 34.175 203.960 34.465 205.125 ;
        RECT 55.650 199.335 57.030 199.505 ;
        RECT 24.480 198.815 24.940 198.985 ;
        RECT 25.740 198.815 27.120 198.985 ;
        RECT 24.565 197.650 24.855 198.815 ;
        RECT 26.080 197.675 26.290 198.815 ;
        RECT 55.990 198.195 56.200 199.335 ;
        RECT 58.190 199.325 58.650 199.495 ;
        RECT 56.370 198.185 56.700 199.165 ;
        RECT 56.470 197.815 56.700 198.185 ;
        RECT 58.275 198.160 58.565 199.325 ;
        RECT 56.470 197.585 57.865 197.815 ;
        RECT 56.370 196.955 56.700 197.585 ;
        RECT 46.490 191.825 48.790 191.995 ;
        RECT 49.720 191.845 50.180 192.015 ;
        RECT 47.005 191.425 47.940 191.825 ;
        RECT 46.575 190.895 47.035 190.915 ;
        RECT 45.370 190.435 47.035 190.895 ;
        RECT 49.805 190.680 50.095 191.845 ;
        RECT 45.370 190.170 46.230 190.435 ;
        RECT 46.575 190.185 47.035 190.435 ;
      LAYER mcon ;
        RECT 31.245 215.735 31.415 215.905 ;
        RECT 31.705 215.735 31.875 215.905 ;
        RECT 32.165 215.735 32.335 215.905 ;
        RECT 23.585 214.725 23.755 214.895 ;
        RECT 25.445 214.715 25.615 214.885 ;
        RECT 25.905 214.715 26.075 214.885 ;
        RECT 26.365 214.715 26.535 214.885 ;
        RECT 33.620 215.725 33.790 215.895 ;
        RECT 24.235 210.425 24.405 210.595 ;
        RECT 25.585 210.425 25.755 210.595 ;
        RECT 26.045 210.425 26.215 210.595 ;
        RECT 26.505 210.425 26.675 210.595 ;
        RECT 41.485 210.025 41.655 210.195 ;
        RECT 41.945 210.025 42.115 210.195 ;
        RECT 42.405 210.025 42.575 210.195 ;
        RECT 42.865 210.025 43.035 210.195 ;
        RECT 43.325 210.025 43.495 210.195 ;
        RECT 43.785 210.025 43.955 210.195 ;
        RECT 44.245 210.025 44.415 210.195 ;
        RECT 45.835 210.025 46.005 210.195 ;
        RECT 53.085 209.975 53.255 210.145 ;
        RECT 53.545 209.975 53.715 210.145 ;
        RECT 54.005 209.975 54.175 210.145 ;
        RECT 54.465 209.975 54.635 210.145 ;
        RECT 54.925 209.975 55.095 210.145 ;
        RECT 56.635 209.975 56.805 210.145 ;
        RECT 24.295 205.055 24.465 205.225 ;
        RECT 25.705 205.075 25.875 205.245 ;
        RECT 26.165 205.075 26.335 205.245 ;
        RECT 26.625 205.075 26.795 205.245 ;
        RECT 31.595 205.105 31.765 205.275 ;
        RECT 32.055 205.105 32.225 205.275 ;
        RECT 32.515 205.105 32.685 205.275 ;
        RECT 34.235 205.125 34.405 205.295 ;
        RECT 55.795 199.335 55.965 199.505 ;
        RECT 56.255 199.335 56.425 199.505 ;
        RECT 56.715 199.335 56.885 199.505 ;
        RECT 24.625 198.815 24.795 198.985 ;
        RECT 25.885 198.815 26.055 198.985 ;
        RECT 26.345 198.815 26.515 198.985 ;
        RECT 26.805 198.815 26.975 198.985 ;
        RECT 58.335 199.325 58.505 199.495 ;
        RECT 57.665 197.615 57.835 197.785 ;
        RECT 46.635 191.825 46.805 191.995 ;
        RECT 47.095 191.825 47.265 191.995 ;
        RECT 47.555 191.825 47.725 191.995 ;
        RECT 48.015 191.825 48.185 191.995 ;
        RECT 48.475 191.825 48.645 191.995 ;
        RECT 49.865 191.845 50.035 192.015 ;
        RECT 45.665 190.465 45.835 190.635 ;
      LAYER met1 ;
        RECT 52.060 217.610 52.565 218.580 ;
        RECT 22.265 215.745 23.785 216.220 ;
        RECT 23.060 215.730 23.785 215.745 ;
        RECT 23.310 215.050 23.785 215.730 ;
        RECT 23.310 215.015 23.900 215.050 ;
        RECT 26.320 215.040 26.780 217.430 ;
        RECT 31.825 216.495 32.320 217.505 ;
        RECT 31.840 216.060 32.300 216.495 ;
        RECT 34.200 216.420 34.700 217.510 ;
        RECT 31.100 215.580 32.480 216.060 ;
        RECT 33.470 215.960 34.700 216.420 ;
        RECT 33.475 215.570 33.935 215.960 ;
        RECT 23.440 214.570 23.900 215.015 ;
        RECT 25.300 214.990 26.780 215.040 ;
        RECT 25.300 214.560 26.680 214.990 ;
        RECT 52.080 212.970 52.540 217.610 ;
        RECT 46.980 212.580 48.040 212.595 ;
        RECT 42.930 212.120 48.040 212.580 ;
        RECT 52.080 212.510 53.970 212.970 ;
        RECT 57.430 212.840 57.915 214.000 ;
        RECT 27.755 211.190 28.965 211.205 ;
        RECT 21.860 210.750 24.530 210.990 ;
        RECT 25.940 210.750 28.965 211.190 ;
        RECT 21.860 210.530 24.550 210.750 ;
        RECT 24.090 210.270 24.550 210.530 ;
        RECT 25.440 210.730 28.965 210.750 ;
        RECT 25.440 210.270 26.820 210.730 ;
        RECT 27.755 210.715 28.965 210.730 ;
        RECT 42.930 210.350 43.390 212.120 ;
        RECT 46.980 212.110 48.040 212.120 ;
        RECT 47.435 210.420 47.940 210.900 ;
        RECT 46.100 210.350 47.940 210.420 ;
        RECT 41.340 209.870 44.560 210.350 ;
        RECT 45.690 209.915 47.940 210.350 ;
        RECT 53.510 210.300 53.970 212.510 ;
        RECT 57.440 210.680 57.900 212.840 ;
        RECT 45.690 209.870 46.150 209.915 ;
        RECT 52.940 209.820 55.240 210.300 ;
        RECT 56.470 210.220 57.900 210.680 ;
        RECT 56.490 209.820 56.950 210.220 ;
        RECT 26.250 206.180 26.710 206.700 ;
        RECT 21.070 205.985 22.420 206.020 ;
        RECT 21.070 205.500 24.590 205.985 ;
        RECT 21.070 205.460 22.420 205.500 ;
        RECT 24.105 205.380 24.590 205.500 ;
        RECT 26.335 205.415 26.625 206.180 ;
        RECT 36.035 205.510 37.085 205.520 ;
        RECT 32.770 205.430 37.085 205.510 ;
        RECT 26.175 205.400 26.625 205.415 ;
        RECT 24.105 205.210 24.610 205.380 ;
        RECT 24.150 204.900 24.610 205.210 ;
        RECT 25.560 204.920 26.940 205.400 ;
        RECT 31.450 205.050 37.085 205.430 ;
        RECT 31.450 204.950 32.830 205.050 ;
        RECT 34.090 204.970 34.550 205.050 ;
        RECT 36.035 205.045 37.085 205.050 ;
        RECT 23.255 200.410 23.850 200.445 ;
        RECT 23.225 199.815 23.880 200.410 ;
        RECT 26.130 200.070 26.655 201.420 ;
        RECT 56.090 200.860 56.590 201.840 ;
        RECT 58.790 201.825 59.305 201.875 ;
        RECT 23.255 199.570 23.850 199.815 ;
        RECT 23.250 199.110 24.950 199.570 ;
        RECT 26.160 199.155 26.620 200.070 ;
        RECT 56.110 199.660 56.570 200.860 ;
        RECT 58.790 200.855 59.320 201.825 ;
        RECT 58.790 200.840 59.305 200.855 ;
        RECT 58.830 200.665 59.290 200.840 ;
        RECT 57.635 200.435 61.535 200.665 ;
        RECT 55.650 199.180 57.030 199.660 ;
        RECT 26.075 199.140 26.620 199.155 ;
        RECT 23.320 199.100 23.780 199.110 ;
        RECT 24.480 198.660 24.940 199.110 ;
        RECT 25.740 198.660 27.120 199.140 ;
        RECT 57.635 197.845 57.865 200.435 ;
        RECT 58.830 200.080 59.290 200.435 ;
        RECT 58.170 199.620 59.290 200.080 ;
        RECT 58.190 199.170 58.650 199.620 ;
        RECT 58.830 199.600 59.290 199.620 ;
        RECT 57.605 197.555 57.895 197.845 ;
        RECT 57.635 197.485 57.865 197.555 ;
        RECT 61.335 195.215 61.565 200.435 ;
        RECT 44.585 195.085 61.565 195.215 ;
        RECT 44.565 194.985 61.565 195.085 ;
        RECT 44.565 194.315 44.840 194.985 ;
        RECT 44.550 193.095 44.845 193.110 ;
        RECT 44.550 192.455 44.850 193.095 ;
        RECT 46.920 193.020 47.415 193.035 ;
        RECT 44.555 192.205 44.850 192.455 ;
        RECT 44.585 190.665 44.815 192.205 ;
        RECT 46.810 192.150 47.415 193.020 ;
        RECT 49.755 192.170 50.175 192.890 ;
        RECT 46.490 191.670 48.790 192.150 ;
        RECT 49.720 191.690 50.180 192.170 ;
        RECT 45.035 190.665 46.065 190.815 ;
        RECT 44.585 190.435 46.065 190.665 ;
        RECT 45.035 190.285 46.065 190.435 ;
      LAYER via ;
        RECT 52.170 218.190 52.430 218.450 ;
        RECT 26.420 217.000 26.680 217.260 ;
        RECT 22.520 215.850 22.780 216.110 ;
        RECT 31.940 217.070 32.200 217.330 ;
        RECT 34.320 217.020 34.580 217.280 ;
        RECT 57.540 213.460 57.800 213.720 ;
        RECT 47.550 212.220 47.810 212.480 ;
        RECT 22.000 210.630 22.260 210.890 ;
        RECT 28.330 210.830 28.590 211.090 ;
        RECT 47.550 210.490 47.810 210.750 ;
        RECT 26.350 206.310 26.610 206.570 ;
        RECT 21.490 205.560 21.750 205.820 ;
        RECT 36.600 205.150 36.860 205.410 ;
        RECT 56.210 201.440 56.470 201.700 ;
        RECT 26.260 200.880 26.520 201.140 ;
        RECT 23.260 199.820 23.840 200.400 ;
        RECT 58.930 201.440 59.190 201.700 ;
        RECT 44.570 194.370 44.830 194.630 ;
        RECT 44.570 192.570 44.830 192.830 ;
        RECT 47.020 192.610 47.280 192.870 ;
        RECT 49.830 192.580 50.110 192.840 ;
      LAYER met2 ;
        RECT 7.905 218.550 8.960 218.570 ;
        RECT 51.820 218.550 53.110 218.570 ;
        RECT 7.905 218.090 57.840 218.550 ;
        RECT 7.905 218.075 8.960 218.090 ;
        RECT 20.010 210.990 20.470 218.090 ;
        RECT 22.420 216.680 22.880 218.090 ;
        RECT 26.320 216.730 26.780 218.090 ;
        RECT 22.415 215.635 22.890 216.680 ;
        RECT 28.230 211.675 28.690 218.090 ;
        RECT 31.840 217.900 32.300 218.090 ;
        RECT 31.830 216.850 32.310 217.900 ;
        RECT 34.220 216.800 34.680 218.090 ;
        RECT 21.425 210.990 22.525 211.005 ;
        RECT 20.010 210.530 22.525 210.990 ;
        RECT 28.210 210.610 28.715 211.675 ;
        RECT 21.390 210.515 22.525 210.530 ;
        RECT 21.390 207.020 21.850 210.515 ;
        RECT 21.390 206.670 26.670 207.020 ;
        RECT 21.390 206.560 26.740 206.670 ;
        RECT 21.390 202.020 21.850 206.560 ;
        RECT 26.210 206.210 26.740 206.560 ;
        RECT 36.500 205.985 36.960 218.090 ;
        RECT 47.450 211.325 47.910 218.090 ;
        RECT 51.820 218.070 53.110 218.090 ;
        RECT 57.440 217.470 57.840 218.090 ;
        RECT 57.440 214.990 57.900 217.470 ;
        RECT 57.440 214.530 60.430 214.990 ;
        RECT 57.440 213.200 57.900 214.530 ;
        RECT 47.435 210.305 47.925 211.325 ;
        RECT 36.490 204.960 36.975 205.985 ;
        RECT 59.970 202.650 60.430 214.530 ;
        RECT 59.970 202.190 64.430 202.650 ;
        RECT 21.390 201.725 26.620 202.020 ;
        RECT 59.970 201.800 60.430 202.190 ;
        RECT 21.390 201.560 26.645 201.725 ;
        RECT 23.320 200.805 23.780 201.560 ;
        RECT 23.290 200.440 23.815 200.805 ;
        RECT 26.140 200.660 26.645 201.560 ;
        RECT 55.990 201.340 60.430 201.800 ;
        RECT 23.255 199.785 23.850 200.440 ;
        RECT 44.570 194.120 44.830 194.780 ;
        RECT 44.585 193.100 44.815 194.120 ;
        RECT 44.555 192.400 44.855 193.100 ;
        RECT 46.825 192.970 47.850 192.980 ;
        RECT 63.970 192.970 64.430 202.190 ;
        RECT 46.660 192.510 64.430 192.970 ;
        RECT 46.825 192.505 47.850 192.510 ;
      LAYER via2 ;
        RECT 8.110 218.180 8.390 218.460 ;
      LAYER met3 ;
        RECT 7.995 218.550 8.505 218.575 ;
        RECT 2.635 218.090 8.505 218.550 ;
        RECT 7.995 218.065 8.505 218.090 ;
      LAYER via3 ;
        RECT 2.705 218.160 3.025 218.480 ;
      LAYER met4 ;
        RECT 1.000 218.550 3.000 220.760 ;
        RECT 1.000 218.090 3.095 218.550 ;
        RECT 1.000 5.000 3.000 218.090 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 33.620 213.410 33.790 213.935 ;
        RECT 23.585 212.410 23.755 212.935 ;
        RECT 24.235 208.110 24.405 208.635 ;
        RECT 45.835 207.710 46.005 208.235 ;
        RECT 56.635 207.660 56.805 208.185 ;
        RECT 24.295 202.740 24.465 203.265 ;
        RECT 34.235 202.810 34.405 203.335 ;
        RECT 24.625 196.500 24.795 197.025 ;
        RECT 58.335 197.010 58.505 197.535 ;
        RECT 49.865 189.530 50.035 190.055 ;
      LAYER li1 ;
        RECT 31.205 213.185 31.445 213.995 ;
        RECT 32.115 213.185 32.385 213.995 ;
        RECT 31.100 213.015 32.480 213.185 ;
        RECT 33.560 213.175 33.850 213.900 ;
        RECT 33.475 213.005 33.935 213.175 ;
        RECT 23.525 212.175 23.815 212.900 ;
        RECT 23.440 212.005 23.900 212.175 ;
        RECT 25.620 212.165 25.850 212.985 ;
        RECT 25.300 211.995 26.680 212.165 ;
        RECT 24.775 209.105 25.025 209.110 ;
        RECT 24.775 208.865 26.090 209.105 ;
        RECT 54.915 208.870 55.155 209.295 ;
        RECT 24.775 208.860 25.025 208.865 ;
        RECT 24.175 207.875 24.465 208.600 ;
        RECT 25.760 207.875 25.990 208.695 ;
        RECT 42.180 208.465 42.730 208.665 ;
        RECT 54.915 208.630 55.920 208.870 ;
        RECT 54.915 208.315 55.155 208.630 ;
        RECT 24.090 207.705 24.550 207.875 ;
        RECT 25.440 207.705 26.820 207.875 ;
        RECT 41.475 207.475 41.805 207.865 ;
        RECT 42.315 207.475 42.645 207.865 ;
        RECT 44.185 207.475 44.475 208.310 ;
        RECT 45.775 207.475 46.065 208.200 ;
        RECT 41.340 207.305 44.560 207.475 ;
        RECT 45.690 207.305 46.150 207.475 ;
        RECT 53.455 207.425 54.390 207.825 ;
        RECT 56.575 207.425 56.865 208.150 ;
        RECT 52.940 207.255 55.240 207.425 ;
        RECT 56.490 207.255 56.950 207.425 ;
        RECT 31.545 204.725 31.875 204.920 ;
        RECT 30.625 204.555 31.875 204.725 ;
        RECT 31.545 204.135 31.875 204.555 ;
        RECT 31.545 203.965 32.225 204.135 ;
        RECT 24.895 203.795 25.225 203.800 ;
        RECT 24.820 203.755 25.540 203.795 ;
        RECT 24.820 203.515 26.210 203.755 ;
        RECT 24.820 203.475 25.540 203.515 ;
        RECT 24.895 203.470 25.225 203.475 ;
        RECT 32.055 203.365 32.225 203.965 ;
        RECT 24.235 202.505 24.525 203.230 ;
        RECT 25.880 202.525 26.110 203.345 ;
        RECT 31.555 202.555 31.795 203.365 ;
        RECT 31.965 202.725 32.295 203.365 ;
        RECT 32.465 202.555 32.735 203.365 ;
        RECT 34.175 202.575 34.465 203.300 ;
        RECT 24.150 202.335 24.610 202.505 ;
        RECT 25.560 202.355 26.940 202.525 ;
        RECT 31.450 202.385 32.830 202.555 ;
        RECT 34.090 202.405 34.550 202.575 ;
        RECT 24.565 196.265 24.855 196.990 ;
        RECT 26.060 196.265 26.290 197.085 ;
        RECT 55.970 196.785 56.200 197.605 ;
        RECT 55.650 196.615 57.030 196.785 ;
        RECT 58.275 196.775 58.565 197.500 ;
        RECT 58.190 196.605 58.650 196.775 ;
        RECT 24.480 196.095 24.940 196.265 ;
        RECT 25.740 196.095 27.120 196.265 ;
        RECT 48.110 191.315 48.705 191.655 ;
        RECT 48.110 189.995 48.285 191.315 ;
        RECT 48.465 190.720 48.705 191.145 ;
        RECT 48.465 190.480 49.350 190.720 ;
        RECT 48.465 190.165 48.705 190.480 ;
        RECT 48.110 189.825 48.705 189.995 ;
        RECT 47.005 189.275 47.940 189.675 ;
        RECT 48.110 189.655 49.485 189.825 ;
        RECT 48.110 189.445 48.705 189.655 ;
        RECT 49.805 189.295 50.095 190.020 ;
        RECT 46.490 189.105 48.790 189.275 ;
        RECT 49.720 189.125 50.180 189.295 ;
      LAYER mcon ;
        RECT 31.245 213.015 31.415 213.185 ;
        RECT 31.705 213.015 31.875 213.185 ;
        RECT 32.165 213.015 32.335 213.185 ;
        RECT 33.620 213.005 33.790 213.175 ;
        RECT 23.585 212.005 23.755 212.175 ;
        RECT 25.445 211.995 25.615 212.165 ;
        RECT 25.905 211.995 26.075 212.165 ;
        RECT 26.365 211.995 26.535 212.165 ;
        RECT 24.815 208.900 24.985 209.070 ;
        RECT 42.365 208.465 42.535 208.635 ;
        RECT 55.715 208.660 55.885 208.830 ;
        RECT 24.235 207.705 24.405 207.875 ;
        RECT 25.585 207.705 25.755 207.875 ;
        RECT 26.045 207.705 26.215 207.875 ;
        RECT 26.505 207.705 26.675 207.875 ;
        RECT 41.485 207.305 41.655 207.475 ;
        RECT 41.945 207.305 42.115 207.475 ;
        RECT 42.405 207.305 42.575 207.475 ;
        RECT 42.865 207.305 43.035 207.475 ;
        RECT 43.325 207.305 43.495 207.475 ;
        RECT 43.785 207.305 43.955 207.475 ;
        RECT 44.245 207.305 44.415 207.475 ;
        RECT 45.835 207.305 46.005 207.475 ;
        RECT 53.085 207.255 53.255 207.425 ;
        RECT 53.545 207.255 53.715 207.425 ;
        RECT 54.005 207.255 54.175 207.425 ;
        RECT 54.465 207.255 54.635 207.425 ;
        RECT 54.925 207.255 55.095 207.425 ;
        RECT 56.635 207.255 56.805 207.425 ;
        RECT 24.975 203.550 25.145 203.720 ;
        RECT 24.295 202.335 24.465 202.505 ;
        RECT 25.705 202.355 25.875 202.525 ;
        RECT 26.165 202.355 26.335 202.525 ;
        RECT 26.625 202.355 26.795 202.525 ;
        RECT 31.595 202.385 31.765 202.555 ;
        RECT 32.055 202.385 32.225 202.555 ;
        RECT 32.515 202.385 32.685 202.555 ;
        RECT 34.235 202.405 34.405 202.575 ;
        RECT 55.795 196.615 55.965 196.785 ;
        RECT 56.255 196.615 56.425 196.785 ;
        RECT 56.715 196.615 56.885 196.785 ;
        RECT 58.335 196.605 58.505 196.775 ;
        RECT 24.625 196.095 24.795 196.265 ;
        RECT 25.885 196.095 26.055 196.265 ;
        RECT 26.345 196.095 26.515 196.265 ;
        RECT 26.805 196.095 26.975 196.265 ;
        RECT 49.095 190.515 49.265 190.685 ;
        RECT 49.315 189.655 49.485 189.825 ;
        RECT 46.635 189.105 46.805 189.275 ;
        RECT 47.095 189.105 47.265 189.275 ;
        RECT 47.555 189.105 47.725 189.275 ;
        RECT 48.015 189.105 48.185 189.275 ;
        RECT 48.475 189.105 48.645 189.275 ;
        RECT 49.865 189.125 50.035 189.295 ;
      LAYER met1 ;
        RECT 31.100 212.955 32.480 213.340 ;
        RECT 33.475 212.955 33.935 213.330 ;
        RECT 31.100 212.860 33.935 212.955 ;
        RECT 31.270 212.850 33.935 212.860 ;
        RECT 31.270 212.800 33.925 212.850 ;
        RECT 8.145 211.995 8.465 212.050 ;
        RECT 23.440 211.995 23.900 212.330 ;
        RECT 25.300 211.995 26.680 212.320 ;
        RECT 8.145 211.840 26.680 211.995 ;
        RECT 8.145 211.790 8.465 211.840 ;
        RECT 20.815 211.255 25.025 211.505 ;
        RECT 13.040 210.425 13.910 210.460 ;
        RECT 20.815 210.425 21.065 211.255 ;
        RECT 24.775 210.970 25.025 211.255 ;
        RECT 13.040 210.175 21.075 210.425 ;
        RECT 13.040 210.140 13.910 210.175 ;
        RECT 24.775 209.170 25.285 210.970 ;
        RECT 24.745 208.800 25.285 209.170 ;
        RECT 24.090 207.625 24.550 208.030 ;
        RECT 24.075 207.550 24.550 207.625 ;
        RECT 24.075 207.465 24.325 207.550 ;
        RECT 9.460 207.310 24.325 207.465 ;
        RECT 9.460 207.140 17.400 207.310 ;
        RECT 24.880 207.140 25.285 208.800 ;
        RECT 25.440 207.550 26.820 208.030 ;
        RECT 25.615 207.140 25.770 207.550 ;
        RECT 31.270 207.140 31.425 212.800 ;
        RECT 42.315 208.365 42.635 208.735 ;
        RECT 55.630 208.625 56.225 208.870 ;
        RECT 9.475 206.985 31.425 207.140 ;
        RECT 39.665 207.985 39.835 208.000 ;
        RECT 42.365 207.985 42.535 208.365 ;
        RECT 39.665 207.815 42.535 207.985 ;
        RECT 10.450 206.965 17.400 206.985 ;
        RECT 13.110 203.660 13.495 204.345 ;
        RECT 13.165 203.565 13.435 203.660 ;
        RECT 13.215 187.435 13.385 203.565 ;
        RECT 16.900 202.355 17.400 206.965 ;
        RECT 24.880 206.615 25.285 206.985 ;
        RECT 20.430 206.285 25.285 206.615 ;
        RECT 20.430 205.285 20.760 206.285 ;
        RECT 20.430 204.930 20.765 205.285 ;
        RECT 20.425 204.530 20.765 204.930 ;
        RECT 24.880 203.830 25.285 206.285 ;
        RECT 39.665 206.185 39.835 207.815 ;
        RECT 41.340 207.150 44.560 207.630 ;
        RECT 45.690 207.150 46.150 207.630 ;
        RECT 29.985 206.015 39.835 206.185 ;
        RECT 29.985 204.725 30.155 206.015 ;
        RECT 39.665 205.250 39.835 206.015 ;
        RECT 42.985 206.430 43.275 207.150 ;
        RECT 45.825 206.430 45.980 207.150 ;
        RECT 52.940 207.100 55.240 207.580 ;
        RECT 54.635 206.430 54.920 207.100 ;
        RECT 42.985 206.275 54.920 206.430 ;
        RECT 41.950 205.250 42.600 205.400 ;
        RECT 39.650 205.050 42.700 205.250 ;
        RECT 30.595 204.725 30.825 204.785 ;
        RECT 29.985 204.555 30.975 204.725 ;
        RECT 30.595 204.495 30.825 204.555 ;
        RECT 24.865 203.440 25.285 203.830 ;
        RECT 24.880 203.390 25.285 203.440 ;
        RECT 24.150 202.355 24.610 202.660 ;
        RECT 25.560 202.385 26.940 202.680 ;
        RECT 31.450 202.385 32.830 202.710 ;
        RECT 25.560 202.355 32.830 202.385 ;
        RECT 16.900 202.230 32.830 202.355 ;
        RECT 34.090 202.250 34.550 202.730 ;
        RECT 16.900 202.200 26.940 202.230 ;
        RECT 16.900 196.100 17.400 202.200 ;
        RECT 24.150 202.180 24.610 202.200 ;
        RECT 24.480 196.100 24.940 196.420 ;
        RECT 25.740 196.100 27.120 196.420 ;
        RECT 34.240 196.100 34.395 202.250 ;
        RECT 39.650 197.655 39.850 205.050 ;
        RECT 41.950 204.900 42.600 205.050 ;
        RECT 42.985 204.480 43.275 206.275 ;
        RECT 43.590 205.250 43.910 205.280 ;
        RECT 55.980 205.250 56.225 208.625 ;
        RECT 56.490 207.100 56.950 207.580 ;
        RECT 43.590 205.080 56.225 205.250 ;
        RECT 43.590 205.050 56.200 205.080 ;
        RECT 43.590 205.020 43.910 205.050 ;
        RECT 56.625 204.480 56.780 207.100 ;
        RECT 42.985 204.325 56.775 204.480 ;
        RECT 39.600 196.850 39.905 197.655 ;
        RECT 39.650 196.100 39.850 196.850 ;
        RECT 42.985 196.615 43.275 204.325 ;
        RECT 55.650 196.655 57.030 196.940 ;
        RECT 58.190 196.655 58.650 196.930 ;
        RECT 55.650 196.615 58.655 196.655 ;
        RECT 42.985 196.460 58.655 196.615 ;
        RECT 42.985 196.100 43.275 196.460 ;
        RECT 58.190 196.450 58.650 196.460 ;
        RECT 16.900 195.605 43.275 196.100 ;
        RECT 16.900 195.600 43.250 195.605 ;
        RECT 37.575 189.105 37.730 195.600 ;
        RECT 39.650 195.370 39.850 195.600 ;
        RECT 39.630 195.240 39.870 195.370 ;
        RECT 39.610 194.460 39.895 195.240 ;
        RECT 39.650 193.550 39.850 194.460 ;
        RECT 39.650 193.350 49.320 193.550 ;
        RECT 39.650 189.105 39.850 193.350 ;
        RECT 49.110 190.720 49.310 193.350 ;
        RECT 49.030 190.700 49.330 190.720 ;
        RECT 49.030 190.500 49.390 190.700 ;
        RECT 49.030 190.480 49.330 190.500 ;
        RECT 49.280 189.460 49.520 189.890 ;
        RECT 46.490 189.105 48.790 189.430 ;
        RECT 37.575 188.950 48.825 189.105 ;
        RECT 48.275 188.330 48.430 188.950 ;
        RECT 48.570 188.330 48.830 188.410 ;
        RECT 48.275 188.175 48.830 188.330 ;
        RECT 48.570 188.090 48.830 188.175 ;
        RECT 49.315 187.435 49.485 189.460 ;
        RECT 49.720 189.105 50.180 189.450 ;
        RECT 49.720 188.970 50.875 189.105 ;
        RECT 49.945 188.950 50.875 188.970 ;
        RECT 49.800 188.330 50.550 188.400 ;
        RECT 50.720 188.330 50.875 188.950 ;
        RECT 49.800 188.175 50.875 188.330 ;
        RECT 49.800 188.100 50.550 188.175 ;
        RECT 13.215 187.265 49.485 187.435 ;
      LAYER via ;
        RECT 8.175 211.790 8.435 212.050 ;
        RECT 13.170 210.170 13.430 210.430 ;
        RECT 9.670 207.095 9.930 207.355 ;
        RECT 13.170 203.920 13.430 204.180 ;
        RECT 20.470 204.670 20.730 204.930 ;
        RECT 42.170 205.020 42.430 205.280 ;
        RECT 43.620 205.020 43.880 205.280 ;
        RECT 39.620 197.020 39.880 197.280 ;
        RECT 39.625 194.920 39.885 195.180 ;
        RECT 48.570 188.120 48.830 188.380 ;
        RECT 49.975 188.125 50.235 188.385 ;
      LAYER met2 ;
        RECT 7.030 212.050 7.470 212.100 ;
        RECT 8.175 212.050 8.435 212.080 ;
        RECT 7.030 211.800 8.435 212.050 ;
        RECT 7.030 211.750 7.470 211.800 ;
        RECT 8.175 211.760 8.435 211.800 ;
        RECT 13.175 210.515 13.425 210.575 ;
        RECT 13.135 210.170 13.470 210.515 ;
        RECT 8.460 206.985 10.140 207.465 ;
        RECT 13.175 204.925 13.425 210.170 ;
        RECT 42.100 205.250 42.650 205.400 ;
        RECT 43.620 205.250 43.880 205.310 ;
        RECT 42.100 205.050 44.150 205.250 ;
        RECT 20.135 204.940 20.795 204.995 ;
        RECT 20.135 204.925 20.815 204.940 ;
        RECT 13.175 204.920 20.815 204.925 ;
        RECT 13.080 204.675 20.815 204.920 ;
        RECT 42.100 204.900 42.650 205.050 ;
        RECT 43.620 204.990 43.880 205.050 ;
        RECT 13.080 203.780 13.525 204.675 ;
        RECT 20.135 204.605 20.815 204.675 ;
        RECT 13.120 203.770 13.485 203.780 ;
        RECT 39.595 196.895 39.905 197.405 ;
        RECT 39.650 195.475 39.850 196.895 ;
        RECT 39.630 195.445 39.875 195.475 ;
        RECT 39.610 194.710 39.895 195.445 ;
        RECT 48.540 188.355 48.860 188.380 ;
        RECT 49.850 188.355 50.460 188.410 ;
        RECT 48.540 188.145 50.460 188.355 ;
        RECT 48.540 188.120 48.860 188.145 ;
        RECT 49.850 188.110 50.460 188.145 ;
      LAYER via2 ;
        RECT 7.110 211.785 7.390 212.065 ;
        RECT 8.610 207.085 8.890 207.365 ;
      LAYER met3 ;
        RECT 5.945 212.100 6.455 212.150 ;
        RECT 7.050 212.100 7.450 212.125 ;
        RECT 5.945 211.750 7.450 212.100 ;
        RECT 5.945 211.700 6.455 211.750 ;
        RECT 7.050 211.725 7.450 211.750 ;
        RECT 8.485 207.465 9.015 207.490 ;
        RECT 7.210 206.985 9.015 207.465 ;
        RECT 8.485 206.960 9.015 206.985 ;
      LAYER via3 ;
        RECT 6.040 211.765 6.360 212.085 ;
        RECT 7.490 207.065 7.810 207.385 ;
      LAYER met4 ;
        RECT 4.000 212.155 6.000 220.760 ;
        RECT 4.000 211.695 6.430 212.155 ;
        RECT 4.000 207.465 6.000 211.695 ;
        RECT 7.405 207.465 7.895 207.470 ;
        RECT 4.000 206.985 7.895 207.465 ;
        RECT 4.000 5.000 6.000 206.985 ;
        RECT 7.405 206.980 7.895 206.985 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 31.250 213.015 31.420 213.185 ;
        RECT 25.445 211.995 25.615 212.165 ;
        RECT 25.585 207.705 25.755 207.875 ;
        RECT 41.485 207.305 41.655 207.475 ;
        RECT 53.090 207.255 53.260 207.425 ;
        RECT 25.705 202.355 25.875 202.525 ;
        RECT 31.600 202.385 31.770 202.555 ;
        RECT 55.795 196.615 55.965 196.785 ;
        RECT 25.885 196.095 26.055 196.265 ;
        RECT 46.640 189.105 46.810 189.275 ;
      LAYER li1 ;
        RECT 31.195 215.355 31.525 215.550 ;
        RECT 30.465 215.185 31.525 215.355 ;
        RECT 31.195 214.765 31.525 215.185 ;
        RECT 31.195 214.595 31.875 214.765 ;
        RECT 26.020 213.565 26.350 214.545 ;
        RECT 30.075 214.175 31.535 214.425 ;
        RECT 31.705 213.995 31.875 214.595 ;
        RECT 32.045 214.175 33.245 214.425 ;
        RECT 26.120 213.215 26.350 213.565 ;
        RECT 31.615 213.355 31.945 213.995 ;
        RECT 26.120 212.985 27.515 213.215 ;
        RECT 26.120 212.965 26.350 212.985 ;
        RECT 26.020 212.335 26.350 212.965 ;
        RECT 26.160 209.275 26.490 210.255 ;
        RECT 26.260 208.915 26.490 209.275 ;
        RECT 41.425 209.175 41.805 209.855 ;
        RECT 42.735 209.345 43.065 209.855 ;
        RECT 43.575 209.345 43.975 209.855 ;
        RECT 42.735 209.175 43.975 209.345 ;
        RECT 44.155 209.265 44.475 209.855 ;
        RECT 53.025 209.405 53.285 209.805 ;
        RECT 26.260 208.685 27.615 208.915 ;
        RECT 26.260 208.675 26.490 208.685 ;
        RECT 26.160 208.045 26.490 208.675 ;
        RECT 41.425 208.215 41.595 209.175 ;
        RECT 44.155 209.095 45.385 209.265 ;
        RECT 53.025 209.235 54.390 209.405 ;
        RECT 41.765 208.835 43.070 209.005 ;
        RECT 44.155 208.925 44.475 209.095 ;
        RECT 53.025 209.045 53.485 209.065 ;
        RECT 51.520 209.015 53.485 209.045 ;
        RECT 41.765 208.385 42.010 208.835 ;
        RECT 42.900 208.635 43.070 208.835 ;
        RECT 43.845 208.755 44.475 208.925 ;
        RECT 42.900 208.465 43.275 208.635 ;
        RECT 43.445 208.215 43.675 208.715 ;
        RECT 41.425 208.045 43.675 208.215 ;
        RECT 41.975 207.725 42.145 208.045 ;
        RECT 43.845 207.875 44.015 208.755 ;
        RECT 51.500 208.615 53.485 209.015 ;
        RECT 51.520 208.585 53.485 208.615 ;
        RECT 53.025 208.335 53.485 208.585 ;
        RECT 53.655 208.165 54.390 209.235 ;
        RECT 43.060 207.705 44.015 207.875 ;
        RECT 53.025 207.995 54.390 208.165 ;
        RECT 53.025 207.595 53.285 207.995 ;
        RECT 26.280 203.925 26.610 204.905 ;
        RECT 26.380 203.615 26.610 203.925 ;
        RECT 31.535 203.790 31.885 203.795 ;
        RECT 26.380 203.385 28.085 203.615 ;
        RECT 30.600 203.545 31.885 203.790 ;
        RECT 32.395 203.545 33.645 203.795 ;
        RECT 26.380 203.325 26.610 203.385 ;
        RECT 26.280 202.695 26.610 203.325 ;
        RECT 26.460 197.665 26.790 198.645 ;
        RECT 55.180 197.775 56.300 198.015 ;
        RECT 26.560 197.315 26.790 197.665 ;
        RECT 26.560 197.085 28.015 197.315 ;
        RECT 26.560 197.065 26.790 197.085 ;
        RECT 26.460 196.435 26.790 197.065 ;
        RECT 46.575 191.255 46.835 191.655 ;
        RECT 46.575 191.085 47.940 191.255 ;
        RECT 47.205 190.015 47.940 191.085 ;
        RECT 46.575 189.845 47.940 190.015 ;
        RECT 46.575 189.445 46.835 189.845 ;
      LAYER mcon ;
        RECT 30.115 214.215 30.285 214.385 ;
        RECT 32.995 214.215 33.165 214.385 ;
        RECT 27.265 213.015 27.435 213.185 ;
        RECT 27.415 208.715 27.585 208.885 ;
        RECT 45.215 209.095 45.385 209.265 ;
        RECT 41.765 208.815 41.935 208.985 ;
        RECT 51.615 208.730 51.785 208.900 ;
        RECT 27.885 203.415 28.055 203.585 ;
        RECT 30.675 203.580 30.845 203.750 ;
        RECT 33.445 203.585 33.615 203.755 ;
        RECT 55.265 197.810 55.435 197.980 ;
        RECT 27.805 197.115 27.975 197.285 ;
      LAYER met1 ;
        RECT 27.675 217.890 33.205 217.895 ;
        RECT 27.675 217.645 33.240 217.890 ;
        RECT 27.685 213.215 27.915 217.645 ;
        RECT 30.405 215.355 30.695 215.385 ;
        RECT 29.765 215.185 30.695 215.355 ;
        RECT 29.765 215.030 29.935 215.185 ;
        RECT 30.405 215.155 30.695 215.185 ;
        RECT 29.690 214.770 30.010 215.030 ;
        RECT 32.960 214.425 33.240 217.645 ;
        RECT 27.185 212.985 27.915 213.215 ;
        RECT 29.525 214.175 30.355 214.425 ;
        RECT 32.915 214.175 33.275 214.425 ;
        RECT 29.525 208.915 29.775 214.175 ;
        RECT 32.960 214.160 33.240 214.175 ;
        RECT 31.940 212.385 32.260 212.430 ;
        RECT 31.940 212.215 39.935 212.385 ;
        RECT 31.940 212.170 32.260 212.215 ;
        RECT 27.355 208.685 29.775 208.915 ;
        RECT 39.765 208.985 39.935 212.215 ;
        RECT 45.215 211.215 51.035 211.235 ;
        RECT 45.185 211.065 51.035 211.215 ;
        RECT 45.185 209.265 45.420 211.065 ;
        RECT 45.115 209.095 45.420 209.265 ;
        RECT 41.665 208.985 42.035 209.085 ;
        RECT 45.185 209.035 45.420 209.095 ;
        RECT 50.570 209.045 51.035 211.065 ;
        RECT 39.765 208.815 42.035 208.985 ;
        RECT 41.665 208.715 42.035 208.815 ;
        RECT 50.570 208.585 51.980 209.045 ;
        RECT 50.580 207.060 50.820 208.585 ;
        RECT 50.570 206.740 50.830 207.060 ;
        RECT 30.640 203.790 30.885 203.820 ;
        RECT 27.825 203.615 28.115 203.645 ;
        RECT 28.410 203.615 31.020 203.790 ;
        RECT 27.765 203.545 31.020 203.615 ;
        RECT 27.765 203.385 28.645 203.545 ;
        RECT 30.640 203.515 30.885 203.545 ;
        RECT 27.825 203.355 28.115 203.385 ;
        RECT 33.330 203.180 33.670 203.820 ;
        RECT 50.570 203.270 50.830 203.730 ;
        RECT 27.745 197.315 28.035 197.345 ;
        RECT 33.360 197.315 33.640 203.180 ;
        RECT 50.430 202.780 50.920 203.270 ;
        RECT 50.580 198.015 50.820 202.780 ;
        RECT 50.580 197.775 55.520 198.015 ;
        RECT 27.705 197.085 33.635 197.315 ;
        RECT 27.745 197.055 28.035 197.085 ;
      LAYER via ;
        RECT 29.720 214.770 29.980 215.030 ;
        RECT 31.970 212.170 32.230 212.430 ;
        RECT 50.570 206.770 50.830 207.030 ;
        RECT 50.570 203.020 50.830 203.280 ;
      LAYER met2 ;
        RECT 29.720 214.740 29.980 215.060 ;
        RECT 29.765 212.385 29.935 214.740 ;
        RECT 31.970 212.385 32.230 212.460 ;
        RECT 29.765 212.215 32.230 212.385 ;
        RECT 31.970 212.140 32.230 212.215 ;
        RECT 50.540 206.770 50.860 207.030 ;
        RECT 50.580 203.520 50.820 206.770 ;
        RECT 50.430 202.880 50.920 203.520 ;
  END
END tt_um_template
END LIBRARY

