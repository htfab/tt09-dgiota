VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_4
  CLASS BLOCK ;
  FOREIGN tt_um_test_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 53.520 142.525 54.115 142.865 ;
        RECT 53.520 141.205 53.695 142.525 ;
        RECT 53.520 141.100 54.115 141.205 ;
        RECT 53.520 140.800 54.900 141.100 ;
        RECT 53.520 140.655 54.115 140.800 ;
      LAYER mcon ;
        RECT 54.630 140.830 54.870 141.070 ;
      LAYER met1 ;
        RECT 54.570 140.800 119.730 141.100 ;
      LAYER via ;
        RECT 119.400 140.800 119.700 141.100 ;
      LAYER met2 ;
        RECT 119.400 83.300 119.700 141.130 ;
        RECT 119.410 83.265 119.690 83.300 ;
      LAYER via2 ;
        RECT 119.410 83.310 119.690 83.590 ;
      LAYER met3 ;
        RECT 119.385 83.600 119.715 83.615 ;
        RECT 119.385 83.300 148.900 83.600 ;
        RECT 119.385 83.285 119.715 83.300 ;
        RECT 148.600 4.000 148.900 83.300 ;
        RECT 148.600 3.700 152.400 4.000 ;
        RECT 152.100 1.340 152.400 3.700 ;
        RECT 152.090 0.960 152.410 1.340 ;
      LAYER via3 ;
        RECT 152.090 0.990 152.410 1.310 ;
      LAYER met4 ;
        RECT 152.085 1.000 152.415 1.315 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 30.520 159.700 30.850 159.715 ;
        RECT 29.350 159.500 30.850 159.700 ;
        RECT 30.520 159.475 30.850 159.500 ;
      LAYER mcon ;
        RECT 29.365 159.515 29.535 159.685 ;
      LAYER met1 ;
        RECT 24.470 159.700 24.730 159.760 ;
        RECT 17.950 159.500 24.730 159.700 ;
        RECT 17.950 135.500 18.250 159.500 ;
        RECT 24.470 159.440 24.730 159.500 ;
        RECT 26.570 159.700 26.830 159.760 ;
        RECT 29.305 159.700 29.595 159.715 ;
        RECT 26.570 159.500 29.595 159.700 ;
        RECT 26.570 159.440 26.830 159.500 ;
        RECT 29.305 159.485 29.595 159.500 ;
        RECT 17.950 135.200 83.080 135.500 ;
      LAYER via ;
        RECT 24.470 159.470 24.730 159.730 ;
        RECT 26.570 159.470 26.830 159.730 ;
        RECT 82.750 135.200 83.050 135.500 ;
      LAYER met2 ;
        RECT 24.440 159.700 24.760 159.730 ;
        RECT 26.540 159.700 26.860 159.730 ;
        RECT 24.440 159.500 26.860 159.700 ;
        RECT 24.440 159.470 24.760 159.500 ;
        RECT 26.540 159.470 26.860 159.500 ;
        RECT 82.750 78.450 83.050 135.530 ;
        RECT 82.760 78.415 83.040 78.450 ;
      LAYER via2 ;
        RECT 82.760 78.460 83.040 78.740 ;
      LAYER met3 ;
        RECT 82.735 78.750 83.065 78.765 ;
        RECT 82.735 78.450 128.750 78.750 ;
        RECT 82.735 78.435 83.065 78.450 ;
        RECT 128.450 1.950 128.750 78.450 ;
        RECT 128.450 1.650 133.100 1.950 ;
        RECT 132.800 1.340 133.100 1.650 ;
        RECT 132.790 0.960 133.110 1.340 ;
      LAYER via3 ;
        RECT 132.790 0.990 133.110 1.310 ;
      LAYER met4 ;
        RECT 132.785 1.000 133.115 1.315 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 32.020 173.850 32.350 173.865 ;
        RECT 31.000 173.650 32.350 173.850 ;
        RECT 32.020 173.625 32.350 173.650 ;
      LAYER mcon ;
        RECT 31.015 173.665 31.185 173.835 ;
      LAYER met1 ;
        RECT 30.955 173.850 31.245 173.865 ;
        RECT 14.750 173.650 31.245 173.850 ;
        RECT 14.750 131.550 15.050 173.650 ;
        RECT 30.955 173.635 31.245 173.650 ;
        RECT 14.750 131.250 77.780 131.550 ;
      LAYER via ;
        RECT 77.450 131.250 77.750 131.550 ;
      LAYER met2 ;
        RECT 77.450 73.600 77.750 131.580 ;
        RECT 77.460 73.565 77.740 73.600 ;
      LAYER via2 ;
        RECT 77.460 73.610 77.740 73.890 ;
      LAYER met3 ;
        RECT 77.435 73.900 77.765 73.915 ;
        RECT 77.435 73.600 109.900 73.900 ;
        RECT 77.435 73.585 77.765 73.600 ;
        RECT 109.600 3.600 109.900 73.600 ;
        RECT 109.600 3.300 113.750 3.600 ;
        RECT 113.450 1.340 113.750 3.300 ;
        RECT 113.440 0.960 113.760 1.340 ;
      LAYER via3 ;
        RECT 113.440 0.990 113.760 1.310 ;
      LAYER met4 ;
        RECT 113.435 1.000 113.765 1.315 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 31.510 175.450 34.550 175.460 ;
        RECT 31.510 173.855 36.290 175.450 ;
        RECT 34.530 173.845 36.290 173.855 ;
        RECT 39.110 172.160 42.150 172.460 ;
        RECT 39.110 170.855 43.900 172.160 ;
        RECT 42.130 170.555 43.900 170.855 ;
        RECT 31.060 170.150 33.650 170.160 ;
        RECT 31.060 168.555 35.190 170.150 ;
        RECT 33.630 168.545 35.190 168.555 ;
        RECT 50.500 163.800 55.400 163.850 ;
        RECT 50.500 162.245 57.190 163.800 ;
        RECT 55.330 162.195 57.190 162.245 ;
        RECT 32.630 161.310 34.340 161.350 ;
        RECT 30.010 159.745 34.340 161.310 ;
        RECT 30.010 159.705 32.750 159.745 ;
        RECT 39.860 158.800 42.900 158.810 ;
        RECT 39.860 157.205 44.590 158.800 ;
        RECT 42.880 157.195 44.590 157.205 ;
        RECT 30.050 154.845 34.190 156.450 ;
        RECT 37.450 145.350 40.050 145.400 ;
        RECT 27.530 145.160 29.190 145.200 ;
        RECT 23.160 143.595 29.190 145.160 ;
        RECT 37.450 143.795 41.540 145.350 ;
        RECT 39.880 143.745 41.540 143.795 ;
        RECT 23.160 143.555 27.550 143.595 ;
        RECT 51.710 143.300 55.800 143.310 ;
        RECT 51.710 141.705 57.540 143.300 ;
        RECT 55.780 141.695 57.540 141.705 ;
      LAYER li1 ;
        RECT 31.700 175.185 33.080 175.355 ;
        RECT 32.040 174.045 32.250 175.185 ;
        RECT 35.640 175.175 36.100 175.345 ;
        RECT 35.725 174.010 36.015 175.175 ;
        RECT 39.300 172.185 40.680 172.355 ;
        RECT 40.255 171.045 40.585 172.185 ;
        RECT 43.250 171.885 43.710 172.055 ;
        RECT 43.335 170.720 43.625 171.885 ;
        RECT 31.250 169.885 32.630 170.055 ;
        RECT 31.590 168.745 31.800 169.885 ;
        RECT 34.540 169.875 35.000 170.045 ;
        RECT 34.625 168.710 34.915 169.875 ;
        RECT 50.690 163.575 53.910 163.745 ;
        RECT 51.745 162.725 51.915 163.575 ;
        RECT 52.585 163.065 52.755 163.575 ;
        RECT 56.540 163.525 57.000 163.695 ;
        RECT 56.625 162.360 56.915 163.525 ;
        RECT 30.200 161.035 31.580 161.205 ;
        RECT 33.690 161.075 34.150 161.245 ;
        RECT 30.540 159.895 30.750 161.035 ;
        RECT 33.775 159.910 34.065 161.075 ;
        RECT 40.050 158.535 41.430 158.705 ;
        RECT 41.005 157.395 41.335 158.535 ;
        RECT 43.940 158.525 44.400 158.695 ;
        RECT 44.025 157.360 44.315 158.525 ;
        RECT 30.240 156.175 31.620 156.345 ;
        RECT 33.540 156.175 34.000 156.345 ;
        RECT 30.580 155.035 30.790 156.175 ;
        RECT 33.625 155.010 33.915 156.175 ;
        RECT 37.640 145.125 39.020 145.295 ;
        RECT 23.350 144.885 25.650 145.055 ;
        RECT 28.540 144.925 29.000 145.095 ;
        RECT 23.865 144.485 24.800 144.885 ;
        RECT 28.625 143.760 28.915 144.925 ;
        RECT 37.980 143.985 38.190 145.125 ;
        RECT 40.890 145.075 41.350 145.245 ;
        RECT 40.975 143.910 41.265 145.075 ;
        RECT 51.900 143.035 54.200 143.205 ;
        RECT 52.415 142.635 53.350 143.035 ;
        RECT 56.890 143.025 57.350 143.195 ;
        RECT 56.975 141.860 57.265 143.025 ;
      LAYER mcon ;
        RECT 31.845 175.185 32.015 175.355 ;
        RECT 32.305 175.185 32.475 175.355 ;
        RECT 32.765 175.185 32.935 175.355 ;
        RECT 35.785 175.175 35.955 175.345 ;
        RECT 39.445 172.185 39.615 172.355 ;
        RECT 39.905 172.185 40.075 172.355 ;
        RECT 40.365 172.185 40.535 172.355 ;
        RECT 43.395 171.885 43.565 172.055 ;
        RECT 31.395 169.885 31.565 170.055 ;
        RECT 31.855 169.885 32.025 170.055 ;
        RECT 32.315 169.885 32.485 170.055 ;
        RECT 34.685 169.875 34.855 170.045 ;
        RECT 50.835 163.575 51.005 163.745 ;
        RECT 51.295 163.575 51.465 163.745 ;
        RECT 51.755 163.575 51.925 163.745 ;
        RECT 52.215 163.575 52.385 163.745 ;
        RECT 52.675 163.575 52.845 163.745 ;
        RECT 53.135 163.575 53.305 163.745 ;
        RECT 53.595 163.575 53.765 163.745 ;
        RECT 56.685 163.525 56.855 163.695 ;
        RECT 30.345 161.035 30.515 161.205 ;
        RECT 30.805 161.035 30.975 161.205 ;
        RECT 31.265 161.035 31.435 161.205 ;
        RECT 33.835 161.075 34.005 161.245 ;
        RECT 40.195 158.535 40.365 158.705 ;
        RECT 40.655 158.535 40.825 158.705 ;
        RECT 41.115 158.535 41.285 158.705 ;
        RECT 44.085 158.525 44.255 158.695 ;
        RECT 30.385 156.175 30.555 156.345 ;
        RECT 30.845 156.175 31.015 156.345 ;
        RECT 31.305 156.175 31.475 156.345 ;
        RECT 33.685 156.175 33.855 156.345 ;
        RECT 37.785 145.125 37.955 145.295 ;
        RECT 38.245 145.125 38.415 145.295 ;
        RECT 38.705 145.125 38.875 145.295 ;
        RECT 23.495 144.885 23.665 145.055 ;
        RECT 23.955 144.885 24.125 145.055 ;
        RECT 24.415 144.885 24.585 145.055 ;
        RECT 24.875 144.885 25.045 145.055 ;
        RECT 25.335 144.885 25.505 145.055 ;
        RECT 28.685 144.925 28.855 145.095 ;
        RECT 41.035 145.075 41.205 145.245 ;
        RECT 52.045 143.035 52.215 143.205 ;
        RECT 52.505 143.035 52.675 143.205 ;
        RECT 52.965 143.035 53.135 143.205 ;
        RECT 53.425 143.035 53.595 143.205 ;
        RECT 53.885 143.035 54.055 143.205 ;
        RECT 57.035 143.025 57.205 143.195 ;
      LAYER met1 ;
        RECT 32.460 176.395 32.750 176.430 ;
        RECT 32.460 176.070 32.765 176.395 ;
        RECT 32.475 175.510 32.765 176.070 ;
        RECT 31.700 175.030 33.080 175.510 ;
        RECT 35.700 175.500 36.000 176.880 ;
        RECT 35.640 175.020 36.100 175.500 ;
        RECT 43.350 173.300 43.650 173.330 ;
        RECT 43.345 172.970 43.650 173.300 ;
        RECT 39.300 172.400 40.680 172.510 ;
        RECT 41.100 172.400 41.400 172.430 ;
        RECT 39.300 172.100 41.400 172.400 ;
        RECT 43.345 172.210 43.645 172.970 ;
        RECT 39.300 172.030 40.680 172.100 ;
        RECT 41.100 172.070 41.400 172.100 ;
        RECT 43.250 171.730 43.710 172.210 ;
        RECT 29.205 170.655 31.855 170.945 ;
        RECT 24.910 170.195 25.200 170.230 ;
        RECT 29.205 170.195 29.495 170.655 ;
        RECT 31.565 170.210 31.855 170.655 ;
        RECT 24.905 169.905 29.495 170.195 ;
        RECT 24.910 169.870 25.200 169.905 ;
        RECT 31.250 169.730 32.630 170.210 ;
        RECT 34.600 170.200 34.895 170.880 ;
        RECT 34.540 169.720 35.000 170.200 ;
        RECT 55.750 164.895 56.900 164.900 ;
        RECT 52.385 164.605 56.900 164.895 ;
        RECT 52.385 163.900 52.675 164.605 ;
        RECT 54.620 164.600 54.980 164.605 ;
        RECT 55.750 164.595 56.900 164.605 ;
        RECT 50.690 163.420 53.910 163.900 ;
        RECT 56.595 163.850 56.900 164.595 ;
        RECT 56.540 163.370 57.000 163.850 ;
        RECT 30.510 162.345 30.800 162.380 ;
        RECT 30.510 162.020 30.805 162.345 ;
        RECT 34.600 162.145 34.895 162.180 ;
        RECT 30.515 161.360 30.805 162.020 ;
        RECT 33.750 161.850 34.895 162.145 ;
        RECT 33.750 161.400 34.045 161.850 ;
        RECT 34.600 161.820 34.895 161.850 ;
        RECT 30.200 160.880 31.580 161.360 ;
        RECT 33.690 160.920 34.150 161.400 ;
        RECT 44.000 159.900 44.300 159.930 ;
        RECT 40.500 159.895 44.300 159.900 ;
        RECT 40.365 159.600 44.300 159.895 ;
        RECT 40.365 158.860 40.655 159.600 ;
        RECT 40.050 158.380 41.430 158.860 ;
        RECT 44.000 158.850 44.300 159.600 ;
        RECT 43.940 158.370 44.400 158.850 ;
        RECT 34.500 156.800 34.800 156.830 ;
        RECT 29.060 156.500 29.350 156.530 ;
        RECT 33.650 156.500 34.800 156.800 ;
        RECT 29.055 156.210 31.620 156.500 ;
        RECT 29.060 156.170 29.350 156.210 ;
        RECT 30.240 156.020 31.620 156.210 ;
        RECT 33.540 156.020 34.000 156.500 ;
        RECT 34.500 156.470 34.800 156.500 ;
        RECT 38.720 146.400 39.085 146.405 ;
        RECT 38.000 146.395 41.250 146.400 ;
        RECT 37.955 146.095 41.250 146.395 ;
        RECT 28.650 146.000 28.955 146.035 ;
        RECT 28.645 145.995 28.955 146.000 ;
        RECT 24.125 145.705 28.955 145.995 ;
        RECT 24.125 145.210 24.415 145.705 ;
        RECT 28.645 145.670 28.955 145.705 ;
        RECT 28.645 145.250 28.950 145.670 ;
        RECT 37.955 145.450 38.245 146.095 ;
        RECT 23.350 144.730 25.650 145.210 ;
        RECT 28.540 144.770 29.000 145.250 ;
        RECT 37.640 144.970 39.020 145.450 ;
        RECT 40.945 145.400 41.250 146.095 ;
        RECT 40.890 144.920 41.350 145.400 ;
        RECT 53.150 144.345 53.440 144.380 ;
        RECT 53.135 144.020 53.440 144.345 ;
        RECT 53.135 143.360 53.425 144.020 ;
        RECT 51.900 142.880 54.200 143.360 ;
        RECT 56.950 143.350 57.250 144.380 ;
        RECT 56.890 142.870 57.350 143.350 ;
      LAYER via ;
        RECT 35.700 176.550 36.000 176.850 ;
        RECT 32.460 176.100 32.750 176.400 ;
        RECT 43.350 173.000 43.650 173.300 ;
        RECT 41.100 172.100 41.400 172.400 ;
        RECT 24.910 169.900 25.200 170.200 ;
        RECT 34.600 170.550 34.895 170.850 ;
        RECT 54.650 164.600 54.950 164.890 ;
        RECT 30.510 162.050 30.800 162.350 ;
        RECT 34.600 161.850 34.895 162.150 ;
        RECT 44.000 159.600 44.300 159.900 ;
        RECT 34.500 156.500 34.800 156.800 ;
        RECT 29.060 156.200 29.350 156.500 ;
        RECT 38.750 146.100 39.055 146.405 ;
        RECT 28.650 145.700 28.955 146.005 ;
        RECT 53.150 144.050 53.440 144.350 ;
        RECT 56.950 144.050 57.250 144.350 ;
      LAYER met2 ;
        RECT 35.060 176.850 35.340 176.885 ;
        RECT 35.050 176.550 36.030 176.850 ;
        RECT 35.060 176.515 35.340 176.550 ;
        RECT 31.760 176.400 32.040 176.435 ;
        RECT 31.750 176.100 32.780 176.400 ;
        RECT 31.760 176.065 32.040 176.100 ;
        RECT 42.510 173.300 42.790 173.335 ;
        RECT 42.500 173.000 43.680 173.300 ;
        RECT 42.510 172.965 42.790 173.000 ;
        RECT 42.010 172.400 42.290 172.435 ;
        RECT 41.070 172.100 42.290 172.400 ;
        RECT 42.010 172.065 42.290 172.100 ;
        RECT 35.560 170.850 35.840 170.885 ;
        RECT 34.570 170.550 35.850 170.850 ;
        RECT 35.560 170.515 35.840 170.550 ;
        RECT 18.960 170.200 19.240 170.235 ;
        RECT 18.950 169.900 25.230 170.200 ;
        RECT 18.960 169.865 19.240 169.900 ;
        RECT 54.650 165.790 54.950 165.800 ;
        RECT 54.615 165.510 54.985 165.790 ;
        RECT 54.650 164.570 54.950 165.510 ;
        RECT 29.760 162.350 30.040 162.385 ;
        RECT 29.750 162.050 30.830 162.350 ;
        RECT 34.570 162.140 35.950 162.150 ;
        RECT 29.760 162.015 30.040 162.050 ;
        RECT 34.570 161.860 35.985 162.140 ;
        RECT 34.570 161.850 35.950 161.860 ;
        RECT 43.970 159.890 45.200 159.900 ;
        RECT 43.970 159.610 45.235 159.890 ;
        RECT 43.970 159.600 45.200 159.610 ;
        RECT 34.470 156.790 35.650 156.800 ;
        RECT 34.470 156.510 35.685 156.790 ;
        RECT 34.470 156.500 35.650 156.510 ;
        RECT 27.900 156.490 29.380 156.500 ;
        RECT 27.865 156.210 29.380 156.490 ;
        RECT 27.900 156.200 29.380 156.210 ;
        RECT 38.760 147.400 39.040 147.435 ;
        RECT 38.750 146.435 39.050 147.400 ;
        RECT 38.750 146.070 39.055 146.435 ;
        RECT 28.620 146.000 28.985 146.005 ;
        RECT 28.620 145.990 30.000 146.000 ;
        RECT 28.620 145.710 30.035 145.990 ;
        RECT 28.620 145.700 30.000 145.710 ;
        RECT 53.120 144.050 57.280 144.350 ;
      LAYER via2 ;
        RECT 35.060 176.560 35.340 176.840 ;
        RECT 31.760 176.110 32.040 176.390 ;
        RECT 42.510 173.010 42.790 173.290 ;
        RECT 42.010 172.110 42.290 172.390 ;
        RECT 35.560 170.560 35.840 170.840 ;
        RECT 18.960 169.910 19.240 170.190 ;
        RECT 21.060 169.910 21.340 170.190 ;
        RECT 54.660 165.510 54.940 165.790 ;
        RECT 29.760 162.060 30.040 162.340 ;
        RECT 35.660 161.860 35.940 162.140 ;
        RECT 44.910 159.610 45.190 159.890 ;
        RECT 35.360 156.510 35.640 156.790 ;
        RECT 27.910 156.210 28.190 156.490 ;
        RECT 38.760 147.110 39.040 147.390 ;
        RECT 29.710 145.710 29.990 145.990 ;
        RECT 55.860 144.060 56.140 144.340 ;
      LAYER met3 ;
        RECT 31.650 179.100 37.750 179.400 ;
        RECT 31.650 177.750 31.950 179.100 ;
        RECT 30.250 177.450 33.850 177.750 ;
        RECT 30.250 176.400 30.550 177.450 ;
        RECT 33.550 176.850 33.850 177.450 ;
        RECT 35.035 176.850 35.365 176.865 ;
        RECT 33.550 176.550 35.365 176.850 ;
        RECT 35.035 176.535 35.365 176.550 ;
        RECT 31.735 176.400 32.065 176.415 ;
        RECT 21.050 176.100 32.065 176.400 ;
        RECT 2.960 170.200 3.340 170.210 ;
        RECT 6.810 170.200 7.190 170.210 ;
        RECT 2.960 169.900 7.190 170.200 ;
        RECT 2.960 169.890 3.340 169.900 ;
        RECT 6.810 169.890 7.190 169.900 ;
        RECT 12.090 170.200 12.410 170.240 ;
        RECT 21.050 170.215 21.350 176.100 ;
        RECT 31.735 176.085 32.065 176.100 ;
        RECT 37.450 175.050 37.750 179.100 ;
        RECT 37.450 174.750 41.950 175.050 ;
        RECT 37.450 172.200 37.750 174.750 ;
        RECT 41.650 174.500 41.950 174.750 ;
        RECT 41.650 174.200 44.600 174.500 ;
        RECT 41.650 173.300 41.950 174.200 ;
        RECT 42.485 173.300 42.815 173.315 ;
        RECT 41.650 173.000 42.815 173.300 ;
        RECT 42.485 172.985 42.815 173.000 ;
        RECT 36.200 171.900 37.750 172.200 ;
        RECT 41.985 172.400 42.315 172.415 ;
        RECT 44.300 172.400 44.600 174.200 ;
        RECT 41.985 172.100 44.600 172.400 ;
        RECT 41.985 172.085 42.315 172.100 ;
        RECT 35.535 170.850 35.865 170.865 ;
        RECT 36.200 170.850 36.500 171.900 ;
        RECT 35.535 170.550 36.500 170.850 ;
        RECT 35.535 170.535 35.865 170.550 ;
        RECT 18.935 170.200 19.265 170.215 ;
        RECT 12.090 169.900 19.265 170.200 ;
        RECT 12.090 169.860 12.410 169.900 ;
        RECT 16.750 168.500 17.050 169.900 ;
        RECT 18.935 169.885 19.265 169.900 ;
        RECT 21.035 169.885 21.365 170.215 ;
        RECT 16.750 168.200 24.200 168.500 ;
        RECT 23.900 162.350 24.200 168.200 ;
        RECT 42.750 166.850 54.950 167.150 ;
        RECT 42.750 163.200 43.050 166.850 ;
        RECT 54.650 165.815 54.950 166.850 ;
        RECT 54.635 165.485 54.965 165.815 ;
        RECT 28.950 162.900 45.200 163.200 ;
        RECT 28.950 162.350 29.250 162.900 ;
        RECT 29.735 162.350 30.065 162.365 ;
        RECT 23.900 162.050 30.065 162.350 ;
        RECT 35.650 162.165 35.950 162.900 ;
        RECT 27.900 157.400 28.200 162.050 ;
        RECT 29.735 162.035 30.065 162.050 ;
        RECT 35.635 161.835 35.965 162.165 ;
        RECT 44.900 159.915 45.200 162.900 ;
        RECT 44.885 159.585 45.215 159.915 ;
        RECT 30.900 157.550 35.650 157.850 ;
        RECT 30.900 157.400 31.200 157.550 ;
        RECT 26.550 157.100 31.200 157.400 ;
        RECT 26.550 149.150 26.850 157.100 ;
        RECT 27.900 156.515 28.200 157.100 ;
        RECT 35.350 156.815 35.650 157.550 ;
        RECT 27.885 156.185 28.215 156.515 ;
        RECT 35.335 156.485 35.665 156.815 ;
        RECT 31.950 151.100 44.450 151.400 ;
        RECT 31.950 149.150 32.250 151.100 ;
        RECT 26.550 148.850 33.800 149.150 ;
        RECT 26.550 147.200 26.850 148.850 ;
        RECT 33.500 147.400 33.800 148.850 ;
        RECT 38.735 147.400 39.065 147.415 ;
        RECT 26.550 146.900 30.000 147.200 ;
        RECT 33.500 147.100 39.065 147.400 ;
        RECT 38.735 147.085 39.065 147.100 ;
        RECT 29.700 146.015 30.000 146.900 ;
        RECT 44.150 146.750 44.450 151.100 ;
        RECT 44.150 146.450 56.150 146.750 ;
        RECT 29.685 145.685 30.015 146.015 ;
        RECT 55.850 144.365 56.150 146.450 ;
        RECT 55.835 144.035 56.165 144.365 ;
      LAYER via3 ;
        RECT 2.990 169.890 3.310 170.210 ;
        RECT 6.840 169.890 7.160 170.210 ;
        RECT 12.090 169.890 12.410 170.210 ;
      LAYER met4 ;
        RECT 1.000 170.215 3.000 220.760 ;
        RECT 1.000 169.885 3.315 170.215 ;
        RECT 6.835 170.200 7.165 170.215 ;
        RECT 12.085 170.200 12.415 170.215 ;
        RECT 6.835 169.900 12.415 170.200 ;
        RECT 6.835 169.885 7.165 169.900 ;
        RECT 12.085 169.885 12.415 169.900 ;
        RECT 1.000 5.000 3.000 169.885 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 35.785 172.860 35.955 173.385 ;
        RECT 43.395 169.570 43.565 170.095 ;
        RECT 34.685 167.560 34.855 168.085 ;
        RECT 56.685 161.210 56.855 161.735 ;
        RECT 33.835 158.760 34.005 159.285 ;
        RECT 44.085 156.210 44.255 156.735 ;
        RECT 33.685 153.860 33.855 154.385 ;
        RECT 28.685 142.610 28.855 143.135 ;
        RECT 41.035 142.760 41.205 143.285 ;
        RECT 57.035 140.710 57.205 141.235 ;
      LAYER li1 ;
        RECT 32.020 172.635 32.250 173.455 ;
        RECT 31.700 172.465 33.080 172.635 ;
        RECT 35.725 172.625 36.015 173.350 ;
        RECT 35.640 172.455 36.100 172.625 ;
        RECT 39.405 169.635 39.645 170.445 ;
        RECT 40.315 169.635 40.585 170.445 ;
        RECT 39.300 169.465 40.680 169.635 ;
        RECT 43.335 169.335 43.625 170.060 ;
        RECT 43.250 169.165 43.710 169.335 ;
        RECT 31.570 167.335 31.800 168.155 ;
        RECT 31.250 167.165 32.630 167.335 ;
        RECT 34.625 167.325 34.915 168.050 ;
        RECT 34.540 167.155 35.000 167.325 ;
        RECT 50.825 161.025 51.155 161.415 ;
        RECT 51.665 161.025 51.995 161.415 ;
        RECT 53.535 161.025 53.825 161.860 ;
        RECT 50.690 160.855 53.910 161.025 ;
        RECT 56.625 160.975 56.915 161.700 ;
        RECT 56.540 160.805 57.000 160.975 ;
        RECT 30.520 158.485 30.750 159.305 ;
        RECT 33.775 158.525 34.065 159.250 ;
        RECT 30.200 158.315 31.580 158.485 ;
        RECT 33.690 158.355 34.150 158.525 ;
        RECT 40.155 155.985 40.395 156.795 ;
        RECT 41.065 155.985 41.335 156.795 ;
        RECT 40.050 155.815 41.430 155.985 ;
        RECT 44.025 155.975 44.315 156.700 ;
        RECT 43.940 155.805 44.400 155.975 ;
        RECT 30.560 153.625 30.790 154.445 ;
        RECT 33.625 153.625 33.915 154.350 ;
        RECT 30.240 153.455 31.620 153.625 ;
        RECT 33.540 153.455 34.000 153.625 ;
        RECT 23.865 142.335 24.800 142.735 ;
        RECT 28.625 142.375 28.915 143.100 ;
        RECT 37.960 142.575 38.190 143.395 ;
        RECT 37.640 142.405 39.020 142.575 ;
        RECT 40.975 142.525 41.265 143.250 ;
        RECT 23.350 142.165 25.650 142.335 ;
        RECT 28.540 142.205 29.000 142.375 ;
        RECT 40.890 142.355 41.350 142.525 ;
        RECT 52.415 140.485 53.350 140.885 ;
        RECT 51.900 140.315 54.200 140.485 ;
        RECT 56.975 140.475 57.265 141.200 ;
        RECT 56.890 140.305 57.350 140.475 ;
      LAYER mcon ;
        RECT 31.845 172.465 32.015 172.635 ;
        RECT 32.305 172.465 32.475 172.635 ;
        RECT 32.765 172.465 32.935 172.635 ;
        RECT 35.785 172.455 35.955 172.625 ;
        RECT 39.445 169.465 39.615 169.635 ;
        RECT 39.905 169.465 40.075 169.635 ;
        RECT 40.365 169.465 40.535 169.635 ;
        RECT 43.395 169.165 43.565 169.335 ;
        RECT 31.395 167.165 31.565 167.335 ;
        RECT 31.855 167.165 32.025 167.335 ;
        RECT 32.315 167.165 32.485 167.335 ;
        RECT 34.685 167.155 34.855 167.325 ;
        RECT 50.835 160.855 51.005 161.025 ;
        RECT 51.295 160.855 51.465 161.025 ;
        RECT 51.755 160.855 51.925 161.025 ;
        RECT 52.215 160.855 52.385 161.025 ;
        RECT 52.675 160.855 52.845 161.025 ;
        RECT 53.135 160.855 53.305 161.025 ;
        RECT 53.595 160.855 53.765 161.025 ;
        RECT 56.685 160.805 56.855 160.975 ;
        RECT 30.345 158.315 30.515 158.485 ;
        RECT 30.805 158.315 30.975 158.485 ;
        RECT 31.265 158.315 31.435 158.485 ;
        RECT 33.835 158.355 34.005 158.525 ;
        RECT 40.195 155.815 40.365 155.985 ;
        RECT 40.655 155.815 40.825 155.985 ;
        RECT 41.115 155.815 41.285 155.985 ;
        RECT 44.085 155.805 44.255 155.975 ;
        RECT 30.385 153.455 30.555 153.625 ;
        RECT 30.845 153.455 31.015 153.625 ;
        RECT 31.305 153.455 31.475 153.625 ;
        RECT 33.685 153.455 33.855 153.625 ;
        RECT 37.785 142.405 37.955 142.575 ;
        RECT 38.245 142.405 38.415 142.575 ;
        RECT 38.705 142.405 38.875 142.575 ;
        RECT 23.495 142.165 23.665 142.335 ;
        RECT 23.955 142.165 24.125 142.335 ;
        RECT 24.415 142.165 24.585 142.335 ;
        RECT 24.875 142.165 25.045 142.335 ;
        RECT 25.335 142.165 25.505 142.335 ;
        RECT 28.685 142.205 28.855 142.375 ;
        RECT 41.035 142.355 41.205 142.525 ;
        RECT 52.045 140.315 52.215 140.485 ;
        RECT 52.505 140.315 52.675 140.485 ;
        RECT 52.965 140.315 53.135 140.485 ;
        RECT 53.425 140.315 53.595 140.485 ;
        RECT 53.885 140.315 54.055 140.485 ;
        RECT 57.035 140.305 57.205 140.475 ;
      LAYER met1 ;
        RECT 31.700 172.310 33.080 172.790 ;
        RECT 24.860 172.045 25.150 172.080 ;
        RECT 32.015 172.045 32.305 172.310 ;
        RECT 35.640 172.300 36.100 172.780 ;
        RECT 24.855 171.755 32.305 172.045 ;
        RECT 35.750 171.770 36.050 172.300 ;
        RECT 24.860 171.720 25.150 171.755 ;
        RECT 38.660 169.600 38.950 169.630 ;
        RECT 39.300 169.600 40.680 169.790 ;
        RECT 38.655 169.310 40.680 169.600 ;
        RECT 38.660 169.270 38.950 169.310 ;
        RECT 43.250 169.010 43.710 169.490 ;
        RECT 43.300 168.270 43.600 169.010 ;
        RECT 31.250 167.010 32.630 167.490 ;
        RECT 26.660 166.495 26.950 166.530 ;
        RECT 31.565 166.495 31.855 167.010 ;
        RECT 34.540 167.000 35.000 167.480 ;
        RECT 26.655 166.205 31.855 166.495 ;
        RECT 34.595 166.680 34.895 167.000 ;
        RECT 34.595 166.350 34.900 166.680 ;
        RECT 34.600 166.320 34.900 166.350 ;
        RECT 26.660 166.170 26.950 166.205 ;
        RECT 49.760 160.990 50.050 161.030 ;
        RECT 50.690 160.990 53.910 161.180 ;
        RECT 49.755 160.700 53.910 160.990 ;
        RECT 49.760 160.670 50.050 160.700 ;
        RECT 56.540 160.650 57.000 161.130 ;
        RECT 56.600 159.720 56.900 160.650 ;
        RECT 30.200 158.160 31.580 158.640 ;
        RECT 33.690 158.250 34.150 158.680 ;
        RECT 34.600 158.250 34.900 158.280 ;
        RECT 33.690 158.200 34.900 158.250 ;
        RECT 26.560 157.845 26.850 157.880 ;
        RECT 30.515 157.845 30.805 158.160 ;
        RECT 33.745 157.950 34.900 158.200 ;
        RECT 34.600 157.920 34.900 157.950 ;
        RECT 26.555 157.555 30.805 157.845 ;
        RECT 26.560 157.520 26.850 157.555 ;
        RECT 39.260 155.950 39.550 155.980 ;
        RECT 40.050 155.950 41.430 156.140 ;
        RECT 39.255 155.660 41.430 155.950 ;
        RECT 39.260 155.620 39.550 155.660 ;
        RECT 43.940 155.650 44.400 156.130 ;
        RECT 44.045 155.085 44.350 155.650 ;
        RECT 44.045 154.750 44.355 155.085 ;
        RECT 44.050 154.720 44.355 154.750 ;
        RECT 30.240 153.300 31.620 153.780 ;
        RECT 33.540 153.300 34.000 153.780 ;
        RECT 30.555 153.130 30.845 153.300 ;
        RECT 30.555 152.805 30.850 153.130 ;
        RECT 30.560 152.770 30.850 152.805 ;
        RECT 33.600 152.600 33.900 153.300 ;
        RECT 33.570 152.300 33.930 152.600 ;
        RECT 36.860 142.540 37.150 142.580 ;
        RECT 37.640 142.540 39.020 142.730 ;
        RECT 23.350 142.010 25.650 142.490 ;
        RECT 28.540 142.050 29.000 142.530 ;
        RECT 36.855 142.250 39.020 142.540 ;
        RECT 36.860 142.220 37.150 142.250 ;
        RECT 40.890 142.200 41.350 142.680 ;
        RECT 29.450 142.050 29.750 142.080 ;
        RECT 24.125 141.780 24.415 142.010 ;
        RECT 24.110 141.455 24.415 141.780 ;
        RECT 28.600 141.750 29.750 142.050 ;
        RECT 40.950 141.950 41.250 142.200 ;
        RECT 29.450 141.720 29.750 141.750 ;
        RECT 40.955 141.700 41.250 141.950 ;
        RECT 24.110 141.420 24.400 141.455 ;
        RECT 40.920 141.405 41.280 141.700 ;
        RECT 51.210 140.450 51.500 140.480 ;
        RECT 51.900 140.450 54.200 140.640 ;
        RECT 51.205 140.160 54.200 140.450 ;
        RECT 51.210 140.120 51.500 140.160 ;
        RECT 56.890 140.150 57.350 140.630 ;
        RECT 56.950 139.420 57.250 140.150 ;
      LAYER via ;
        RECT 24.860 171.750 25.150 172.050 ;
        RECT 35.750 171.800 36.050 172.100 ;
        RECT 38.660 169.300 38.950 169.600 ;
        RECT 43.300 168.300 43.600 168.600 ;
        RECT 26.660 166.200 26.950 166.500 ;
        RECT 34.600 166.350 34.900 166.650 ;
        RECT 49.760 160.700 50.050 161.000 ;
        RECT 56.600 159.750 56.900 160.050 ;
        RECT 26.560 157.550 26.850 157.850 ;
        RECT 34.600 157.950 34.900 158.250 ;
        RECT 39.260 155.650 39.550 155.950 ;
        RECT 44.050 154.750 44.355 155.055 ;
        RECT 30.560 152.800 30.850 153.100 ;
        RECT 33.600 152.300 33.900 152.600 ;
        RECT 36.860 142.250 37.150 142.550 ;
        RECT 29.450 141.750 29.750 142.050 ;
        RECT 24.110 141.450 24.400 141.750 ;
        RECT 40.950 141.405 41.250 141.700 ;
        RECT 51.210 140.150 51.500 140.450 ;
        RECT 56.950 139.450 57.250 139.750 ;
      LAYER met2 ;
        RECT 18.960 172.050 19.240 172.085 ;
        RECT 18.950 171.750 25.180 172.050 ;
        RECT 32.550 171.800 36.080 172.100 ;
        RECT 18.960 171.715 19.240 171.750 ;
        RECT 32.550 166.650 32.850 171.800 ;
        RECT 36.700 169.300 38.980 169.600 ;
        RECT 36.700 168.600 37.000 169.300 ;
        RECT 36.700 168.300 43.630 168.600 ;
        RECT 20.060 166.500 20.340 166.535 ;
        RECT 20.050 166.200 26.980 166.500 ;
        RECT 32.550 166.350 34.930 166.650 ;
        RECT 20.060 166.165 20.340 166.200 ;
        RECT 22.000 164.300 22.300 166.200 ;
        RECT 32.550 164.300 32.850 166.350 ;
        RECT 36.700 164.300 37.000 168.300 ;
        RECT 22.000 164.000 37.000 164.300 ;
        RECT 22.000 157.850 22.300 164.000 ;
        RECT 36.700 161.000 37.000 164.000 ;
        RECT 36.700 160.700 50.080 161.000 ;
        RECT 36.700 158.250 37.000 160.700 ;
        RECT 48.200 160.050 48.500 160.700 ;
        RECT 48.200 159.750 56.930 160.050 ;
        RECT 34.570 157.950 37.000 158.250 ;
        RECT 22.000 157.550 26.880 157.850 ;
        RECT 22.000 153.100 22.300 157.550 ;
        RECT 36.700 155.950 37.000 157.950 ;
        RECT 36.700 155.650 39.580 155.950 ;
        RECT 38.400 155.050 38.700 155.650 ;
        RECT 44.020 155.050 44.385 155.055 ;
        RECT 38.400 154.750 44.385 155.050 ;
        RECT 22.000 152.800 30.880 153.100 ;
        RECT 22.000 141.750 22.300 152.800 ;
        RECT 29.700 151.750 30.000 152.800 ;
        RECT 33.600 151.750 33.900 152.630 ;
        RECT 29.700 151.450 33.900 151.750 ;
        RECT 32.100 142.250 37.180 142.550 ;
        RECT 32.100 142.050 32.400 142.250 ;
        RECT 29.420 141.750 32.400 142.050 ;
        RECT 22.000 141.450 24.430 141.750 ;
        RECT 22.000 139.500 22.300 141.450 ;
        RECT 32.100 140.450 32.400 141.750 ;
        RECT 40.950 140.450 41.250 141.730 ;
        RECT 32.100 140.150 51.530 140.450 ;
        RECT 32.100 139.500 32.400 140.150 ;
        RECT 22.000 139.200 32.400 139.500 ;
        RECT 50.500 138.950 50.800 140.150 ;
        RECT 55.800 139.450 57.280 139.750 ;
        RECT 55.800 138.950 56.100 139.450 ;
        RECT 50.500 138.650 56.100 138.950 ;
      LAYER via2 ;
        RECT 18.960 171.760 19.240 172.040 ;
        RECT 20.060 166.210 20.340 166.490 ;
      LAYER met3 ;
        RECT 12.060 172.050 12.440 172.060 ;
        RECT 18.935 172.050 19.265 172.065 ;
        RECT 12.060 171.750 19.265 172.050 ;
        RECT 12.060 171.740 12.440 171.750 ;
        RECT 18.935 171.735 19.265 171.750 ;
        RECT 12.210 166.500 12.590 166.510 ;
        RECT 20.035 166.500 20.365 166.515 ;
        RECT 12.210 166.200 20.365 166.500 ;
        RECT 12.210 166.190 12.590 166.200 ;
        RECT 20.035 166.185 20.365 166.200 ;
      LAYER via3 ;
        RECT 12.090 171.740 12.410 172.060 ;
        RECT 12.240 166.190 12.560 166.510 ;
      LAYER met4 ;
        RECT 4.000 172.050 6.000 220.760 ;
        RECT 12.085 172.050 12.415 172.065 ;
        RECT 4.000 171.750 12.415 172.050 ;
        RECT 4.000 166.500 6.000 171.750 ;
        RECT 12.085 171.735 12.415 171.750 ;
        RECT 12.235 166.500 12.565 166.515 ;
        RECT 4.000 166.200 12.565 166.500 ;
        RECT 4.000 5.000 6.000 166.200 ;
        RECT 12.235 166.185 12.565 166.200 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 31.845 172.465 32.015 172.635 ;
        RECT 39.450 169.465 39.620 169.635 ;
        RECT 31.395 167.165 31.565 167.335 ;
        RECT 50.835 160.855 51.005 161.025 ;
        RECT 30.345 158.315 30.515 158.485 ;
        RECT 40.200 155.815 40.370 155.985 ;
        RECT 30.385 153.455 30.555 153.625 ;
        RECT 37.785 142.405 37.955 142.575 ;
        RECT 23.500 142.165 23.670 142.335 ;
        RECT 52.050 140.315 52.220 140.485 ;
      LAYER li1 ;
        RECT 32.420 174.035 32.750 175.015 ;
        RECT 32.520 173.715 32.750 174.035 ;
        RECT 32.520 173.485 34.115 173.715 ;
        RECT 32.520 173.435 32.750 173.485 ;
        RECT 32.420 172.805 32.750 173.435 ;
        RECT 38.650 172.900 39.300 173.100 ;
        RECT 38.650 171.750 38.850 172.900 ;
        RECT 39.395 171.750 39.725 172.000 ;
        RECT 38.650 171.550 39.725 171.750 ;
        RECT 39.395 171.215 39.725 171.550 ;
        RECT 39.395 171.045 40.075 171.215 ;
        RECT 39.385 170.625 39.735 170.875 ;
        RECT 39.905 170.445 40.075 171.045 ;
        RECT 40.245 170.845 40.595 170.875 ;
        RECT 40.245 170.655 41.795 170.845 ;
        RECT 40.245 170.625 40.595 170.655 ;
        RECT 39.815 169.805 40.145 170.445 ;
        RECT 31.970 168.735 32.300 169.715 ;
        RECT 31.570 168.550 31.900 168.565 ;
        RECT 30.450 168.350 31.900 168.550 ;
        RECT 31.570 168.325 31.900 168.350 ;
        RECT 32.070 168.415 32.300 168.735 ;
        RECT 32.070 168.185 33.565 168.415 ;
        RECT 32.070 168.135 32.300 168.185 ;
        RECT 31.970 167.505 32.300 168.135 ;
        RECT 50.775 162.725 51.155 163.405 ;
        RECT 52.085 162.895 52.415 163.405 ;
        RECT 52.925 162.895 53.325 163.405 ;
        RECT 52.085 162.725 53.325 162.895 ;
        RECT 53.505 162.750 53.825 163.405 ;
        RECT 50.775 161.765 50.945 162.725 ;
        RECT 51.115 162.385 52.420 162.555 ;
        RECT 53.505 162.475 53.900 162.750 ;
        RECT 51.115 161.935 51.360 162.385 ;
        RECT 51.530 162.015 52.080 162.215 ;
        RECT 52.250 162.185 52.420 162.385 ;
        RECT 53.195 162.450 53.900 162.475 ;
        RECT 53.195 162.305 53.825 162.450 ;
        RECT 52.250 162.015 52.625 162.185 ;
        RECT 52.795 161.765 53.025 162.265 ;
        RECT 50.775 161.595 53.025 161.765 ;
        RECT 51.325 161.275 51.495 161.595 ;
        RECT 53.195 161.425 53.365 162.305 ;
        RECT 52.410 161.255 53.365 161.425 ;
        RECT 30.920 159.885 31.250 160.865 ;
        RECT 31.020 159.515 31.250 159.885 ;
        RECT 31.020 159.285 32.565 159.515 ;
        RECT 30.920 158.655 31.250 159.285 ;
        RECT 32.335 159.135 32.565 159.285 ;
        RECT 40.145 158.100 40.475 158.350 ;
        RECT 40.000 157.800 40.475 158.100 ;
        RECT 40.145 157.565 40.475 157.800 ;
        RECT 40.145 157.395 40.825 157.565 ;
        RECT 39.075 156.975 40.485 157.225 ;
        RECT 40.655 156.795 40.825 157.395 ;
        RECT 40.995 157.200 41.345 157.225 ;
        RECT 40.995 157.000 42.300 157.200 ;
        RECT 40.995 156.975 41.345 157.000 ;
        RECT 40.565 156.155 40.895 156.795 ;
        RECT 30.960 155.025 31.290 156.005 ;
        RECT 30.560 154.850 30.890 154.855 ;
        RECT 29.400 154.650 30.890 154.850 ;
        RECT 30.560 154.615 30.890 154.650 ;
        RECT 31.060 154.665 31.290 155.025 ;
        RECT 32.335 154.665 32.565 154.915 ;
        RECT 31.060 154.435 32.565 154.665 ;
        RECT 31.060 154.425 31.290 154.435 ;
        RECT 30.960 153.795 31.290 154.425 ;
        RECT 23.435 144.315 23.695 144.715 ;
        RECT 24.970 144.375 25.565 144.715 ;
        RECT 23.435 144.145 24.800 144.315 ;
        RECT 23.435 143.500 23.895 143.975 ;
        RECT 22.600 143.300 23.895 143.500 ;
        RECT 23.435 143.245 23.895 143.300 ;
        RECT 24.065 143.075 24.800 144.145 ;
        RECT 23.435 142.905 24.800 143.075 ;
        RECT 24.970 143.055 25.145 144.375 ;
        RECT 25.325 143.450 25.565 144.205 ;
        RECT 38.360 143.975 38.690 144.955 ;
        RECT 37.960 143.800 38.290 143.805 ;
        RECT 36.850 143.600 38.290 143.800 ;
        RECT 37.960 143.565 38.290 143.600 ;
        RECT 25.325 143.250 26.500 143.450 ;
        RECT 38.460 143.375 38.690 143.975 ;
        RECT 25.325 143.225 25.565 143.250 ;
        RECT 23.435 142.505 23.695 142.905 ;
        RECT 24.970 142.505 25.565 143.055 ;
        RECT 38.360 142.745 38.690 143.375 ;
        RECT 51.985 142.465 52.245 142.865 ;
        RECT 51.985 142.295 53.350 142.465 ;
        RECT 51.985 141.650 52.445 142.125 ;
        RECT 51.100 141.450 52.445 141.650 ;
        RECT 51.985 141.395 52.445 141.450 ;
        RECT 52.615 141.225 53.350 142.295 ;
        RECT 53.875 141.650 54.115 142.355 ;
        RECT 53.875 141.450 55.200 141.650 ;
        RECT 53.875 141.375 54.115 141.450 ;
        RECT 51.985 141.055 53.350 141.225 ;
        RECT 51.985 140.655 52.245 141.055 ;
      LAYER mcon ;
        RECT 33.915 173.515 34.085 173.685 ;
        RECT 39.065 172.915 39.235 173.085 ;
        RECT 39.515 170.665 39.685 170.835 ;
        RECT 41.615 170.665 41.785 170.835 ;
        RECT 30.465 168.365 30.635 168.535 ;
        RECT 53.640 162.500 53.840 162.700 ;
        RECT 51.115 162.075 51.285 162.245 ;
        RECT 51.530 162.045 51.700 162.215 ;
        RECT 32.365 159.215 32.535 159.385 ;
        RECT 40.085 157.850 40.285 158.050 ;
        RECT 39.255 157.005 39.445 157.195 ;
        RECT 42.065 157.015 42.235 157.185 ;
        RECT 29.415 154.665 29.585 154.835 ;
        RECT 32.360 154.610 32.540 154.790 ;
        RECT 22.615 143.315 22.785 143.485 ;
        RECT 38.465 143.515 38.635 143.685 ;
        RECT 26.315 143.265 26.485 143.435 ;
        RECT 25.365 142.715 25.535 142.885 ;
        RECT 51.115 141.465 51.285 141.635 ;
        RECT 55.015 141.465 55.185 141.635 ;
      LAYER met1 ;
        RECT 33.885 178.285 38.365 178.515 ;
        RECT 33.885 173.455 34.115 178.285 ;
        RECT 33.335 171.185 37.365 171.415 ;
        RECT 30.405 168.550 30.695 168.565 ;
        RECT 25.450 168.350 30.695 168.550 ;
        RECT 25.450 154.850 25.650 168.350 ;
        RECT 30.405 168.335 30.695 168.350 ;
        RECT 33.335 168.185 33.565 171.185 ;
        RECT 37.135 168.665 37.365 171.185 ;
        RECT 38.135 170.865 38.365 178.285 ;
        RECT 41.050 173.900 45.600 174.100 ;
        RECT 39.005 173.100 39.295 173.115 ;
        RECT 41.050 173.100 41.250 173.900 ;
        RECT 39.000 172.900 41.250 173.100 ;
        RECT 39.005 172.885 39.295 172.900 ;
        RECT 38.135 170.635 39.745 170.865 ;
        RECT 41.585 168.665 41.815 170.895 ;
        RECT 37.135 168.435 41.815 168.665 ;
        RECT 32.335 162.535 38.665 162.765 ;
        RECT 32.335 159.155 32.565 162.535 ;
        RECT 32.335 157.285 36.815 157.515 ;
        RECT 29.355 154.850 29.645 154.865 ;
        RECT 25.450 154.650 29.645 154.850 ;
        RECT 32.335 154.820 32.565 157.285 ;
        RECT 25.450 149.000 25.650 154.650 ;
        RECT 29.355 154.635 29.645 154.650 ;
        RECT 32.330 154.580 32.570 154.820 ;
        RECT 32.335 154.435 32.565 154.580 ;
        RECT 36.585 154.515 36.815 157.285 ;
        RECT 38.435 157.215 38.665 162.535 ;
        RECT 45.400 162.550 45.600 173.900 ;
        RECT 48.200 166.350 61.050 166.550 ;
        RECT 48.200 162.550 48.400 166.350 ;
        RECT 53.550 162.550 55.300 162.750 ;
        RECT 45.400 162.350 50.050 162.550 ;
        RECT 53.580 162.470 53.900 162.550 ;
        RECT 49.775 162.335 50.050 162.350 ;
        RECT 49.775 162.275 51.275 162.335 ;
        RECT 49.775 162.185 51.345 162.275 ;
        RECT 51.055 162.045 51.345 162.185 ;
        RECT 51.500 162.200 51.730 162.275 ;
        RECT 51.500 162.050 52.075 162.200 ;
        RECT 51.500 161.985 51.730 162.050 ;
        RECT 51.500 161.700 51.700 161.985 ;
        RECT 39.250 161.500 51.700 161.700 ;
        RECT 39.250 158.050 39.450 161.500 ;
        RECT 40.055 158.050 40.315 158.080 ;
        RECT 39.250 157.850 40.400 158.050 ;
        RECT 40.055 157.820 40.315 157.850 ;
        RECT 39.195 157.215 39.505 157.225 ;
        RECT 38.435 156.985 39.505 157.215 ;
        RECT 42.005 156.985 42.965 157.215 ;
        RECT 39.195 156.975 39.505 156.985 ;
        RECT 42.735 154.515 42.965 156.985 ;
        RECT 36.585 154.285 42.965 154.515 ;
        RECT 55.100 150.500 55.300 162.550 ;
        RECT 20.100 148.800 25.650 149.000 ;
        RECT 36.850 150.300 55.300 150.500 ;
        RECT 20.100 140.100 20.300 148.800 ;
        RECT 22.600 146.550 35.150 146.750 ;
        RECT 22.600 143.545 22.800 146.550 ;
        RECT 22.585 143.255 22.815 143.545 ;
        RECT 26.255 143.450 26.545 143.465 ;
        RECT 26.255 143.250 27.750 143.450 ;
        RECT 26.255 143.235 26.545 143.250 ;
        RECT 25.305 142.900 25.595 142.915 ;
        RECT 25.305 142.700 26.800 142.900 ;
        RECT 25.305 142.685 25.595 142.700 ;
        RECT 26.600 140.100 26.800 142.700 ;
        RECT 27.550 141.300 27.750 143.250 ;
        RECT 27.550 141.100 32.400 141.300 ;
        RECT 20.100 139.900 26.800 140.100 ;
        RECT 32.200 139.050 32.400 141.100 ;
        RECT 34.950 141.150 35.150 146.550 ;
        RECT 36.850 143.860 37.050 150.300 ;
        RECT 36.820 143.540 37.080 143.860 ;
        RECT 38.405 143.700 38.695 143.715 ;
        RECT 38.405 143.500 40.350 143.700 ;
        RECT 38.405 143.485 38.695 143.500 ;
        RECT 40.150 141.150 40.350 143.500 ;
        RECT 43.650 142.150 43.850 150.300 ;
        RECT 60.850 148.550 61.050 166.350 ;
        RECT 46.400 148.350 61.050 148.550 ;
        RECT 46.400 145.050 46.600 148.350 ;
        RECT 46.400 144.850 55.200 145.050 ;
        RECT 45.320 142.150 45.580 142.210 ;
        RECT 43.650 141.950 45.580 142.150 ;
        RECT 45.320 141.890 45.580 141.950 ;
        RECT 34.950 140.950 40.350 141.150 ;
        RECT 46.400 139.050 46.600 144.850 ;
        RECT 47.420 142.150 47.680 142.210 ;
        RECT 47.420 141.950 51.300 142.150 ;
        RECT 47.420 141.890 47.680 141.950 ;
        RECT 51.100 141.695 51.300 141.950 ;
        RECT 55.000 141.695 55.200 144.850 ;
        RECT 51.085 141.405 51.315 141.695 ;
        RECT 54.985 141.405 55.215 141.695 ;
        RECT 32.200 138.850 46.600 139.050 ;
      LAYER via ;
        RECT 45.320 141.920 45.580 142.180 ;
        RECT 47.420 141.920 47.680 142.180 ;
      LAYER met2 ;
        RECT 45.290 142.150 45.610 142.180 ;
        RECT 47.390 142.150 47.710 142.180 ;
        RECT 45.290 141.950 47.710 142.150 ;
        RECT 45.290 141.920 45.610 141.950 ;
        RECT 47.390 141.920 47.710 141.950 ;
  END
END tt_um_test_3
END LIBRARY

