VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dgiota
  CLASS BLOCK ;
  FOREIGN dgiota ;
  ORIGIN -1.000 0.000 ;
  SIZE 151.710 BY 225.760 ;
  PIN ua[0]
    ANTENNADIFFAREA 0.601000 ;
    PORT
      LAYER li1 ;
        RECT 63.885 70.895 65.505 71.865 ;
        RECT 63.885 70.225 64.225 70.895 ;
        RECT 63.885 69.655 64.355 70.225 ;
      LAYER mcon ;
        RECT 63.945 70.165 64.115 70.335 ;
      LAYER met1 ;
        RECT 63.870 70.120 64.190 70.380 ;
      LAYER via ;
        RECT 63.900 70.120 64.160 70.380 ;
      LAYER met2 ;
        RECT 63.900 70.090 64.160 70.410 ;
        RECT 63.960 69.925 64.100 70.090 ;
        RECT 63.890 69.555 64.170 69.925 ;
      LAYER via2 ;
        RECT 63.890 69.600 64.170 69.880 ;
      LAYER met3 ;
        RECT 44.400 70.040 45.360 70.190 ;
        RECT 44.400 69.890 52.000 70.040 ;
        RECT 63.865 69.890 64.195 69.905 ;
        RECT 44.400 69.590 64.195 69.890 ;
        RECT 44.400 69.440 52.000 69.590 ;
        RECT 63.865 69.575 64.195 69.590 ;
        RECT 44.400 69.290 45.360 69.440 ;
      LAYER via3 ;
        RECT 44.430 69.290 45.330 70.190 ;
      LAYER met4 ;
        RECT 40.270 111.890 152.710 112.790 ;
        RECT 40.270 70.210 41.170 111.890 ;
        RECT 40.270 69.310 45.360 70.210 ;
        RECT 44.425 69.285 45.335 69.310 ;
        RECT 151.810 0.000 152.710 111.890 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 57.005 64.945 57.345 65.315 ;
      LAYER mcon ;
        RECT 57.045 65.065 57.215 65.235 ;
      LAYER met1 ;
        RECT 56.985 65.220 57.275 65.265 ;
        RECT 63.870 65.220 64.190 65.280 ;
        RECT 56.985 65.080 64.190 65.220 ;
        RECT 56.985 65.035 57.275 65.080 ;
        RECT 63.870 65.020 64.190 65.080 ;
      LAYER via ;
        RECT 63.900 65.020 64.160 65.280 ;
      LAYER met2 ;
        RECT 63.900 64.990 64.160 65.310 ;
        RECT 63.960 63.125 64.100 64.990 ;
        RECT 63.890 62.755 64.170 63.125 ;
      LAYER via2 ;
        RECT 63.890 62.800 64.170 63.080 ;
      LAYER met3 ;
        RECT 44.700 63.240 45.660 63.390 ;
        RECT 44.700 63.090 52.000 63.240 ;
        RECT 63.865 63.090 64.195 63.105 ;
        RECT 44.700 62.790 64.195 63.090 ;
        RECT 44.700 62.640 52.000 62.790 ;
        RECT 63.865 62.775 64.195 62.790 ;
        RECT 44.700 62.490 45.660 62.640 ;
      LAYER via3 ;
        RECT 44.730 62.490 45.630 63.390 ;
      LAYER met4 ;
        RECT 44.725 63.390 45.635 63.395 ;
        RECT 40.140 62.490 45.635 63.390 ;
        RECT 40.140 18.330 41.040 62.490 ;
        RECT 44.725 62.485 45.635 62.490 ;
        RECT 40.140 17.430 133.390 18.330 ;
        RECT 132.490 0.000 133.390 17.430 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 57.005 68.045 57.345 68.415 ;
      LAYER mcon ;
        RECT 57.045 68.125 57.215 68.295 ;
      LAYER met1 ;
        RECT 53.750 68.280 54.070 68.340 ;
        RECT 56.985 68.280 57.275 68.325 ;
        RECT 53.750 68.140 57.275 68.280 ;
        RECT 53.750 68.080 54.070 68.140 ;
        RECT 56.985 68.095 57.275 68.140 ;
      LAYER via ;
        RECT 53.780 68.080 54.040 68.340 ;
      LAYER met2 ;
        RECT 53.780 68.050 54.040 68.370 ;
        RECT 53.840 66.525 53.980 68.050 ;
        RECT 53.770 66.155 54.050 66.525 ;
      LAYER via2 ;
        RECT 53.770 66.200 54.050 66.480 ;
      LAYER met3 ;
        RECT 44.715 66.640 45.685 66.795 ;
        RECT 44.715 66.490 52.000 66.640 ;
        RECT 53.745 66.490 54.075 66.505 ;
        RECT 44.715 66.190 54.075 66.490 ;
        RECT 44.715 66.040 52.000 66.190 ;
        RECT 53.745 66.175 54.075 66.190 ;
        RECT 44.715 65.885 45.685 66.040 ;
      LAYER via3 ;
        RECT 44.745 65.885 45.655 66.795 ;
      LAYER met4 ;
        RECT 37.635 66.800 45.545 66.835 ;
        RECT 37.635 65.925 45.660 66.800 ;
        RECT 37.635 14.910 38.545 65.925 ;
        RECT 44.740 65.880 45.660 65.925 ;
        RECT 37.635 14.010 114.070 14.910 ;
        RECT 37.635 14.005 38.545 14.010 ;
        RECT 113.170 0.000 114.070 14.010 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN VDPWR
    ANTENNAGATEAREA 1069.782959 ;
    ANTENNADIFFAREA 255.487289 ;
    PORT
      LAYER nwell ;
        RECT 55.330 97.905 144.490 100.735 ;
        RECT 55.330 92.465 144.490 95.295 ;
        RECT 55.330 87.025 144.490 89.855 ;
        RECT 55.330 81.585 144.490 84.415 ;
        RECT 55.330 76.145 144.490 78.975 ;
        RECT 55.330 70.705 144.490 73.535 ;
        RECT 55.330 65.265 144.490 68.095 ;
        RECT 55.330 59.825 144.490 62.655 ;
        RECT 55.330 54.385 144.490 57.215 ;
        RECT 55.330 48.945 144.490 51.775 ;
        RECT 55.330 43.505 144.490 46.335 ;
        RECT 55.330 38.065 144.490 40.895 ;
        RECT 55.330 32.625 144.490 35.455 ;
        RECT 55.330 27.185 144.490 30.015 ;
      LAYER li1 ;
        RECT 56.295 100.495 56.815 101.035 ;
        RECT 55.605 99.405 56.815 100.495 ;
        RECT 60.390 99.840 60.740 101.090 ;
        RECT 65.910 99.840 66.260 101.090 ;
        RECT 56.985 99.405 62.330 99.840 ;
        RECT 62.505 99.405 67.850 99.840 ;
        RECT 68.485 99.405 68.775 100.570 ;
        RECT 72.350 99.840 72.700 101.090 ;
        RECT 77.870 99.840 78.220 101.090 ;
        RECT 80.675 100.495 81.195 101.035 ;
        RECT 68.945 99.405 74.290 99.840 ;
        RECT 74.465 99.405 79.810 99.840 ;
        RECT 79.985 99.405 81.195 100.495 ;
        RECT 81.365 99.405 81.655 100.570 ;
        RECT 85.230 99.840 85.580 101.090 ;
        RECT 90.750 99.840 91.100 101.090 ;
        RECT 93.555 100.495 94.075 101.035 ;
        RECT 81.825 99.405 87.170 99.840 ;
        RECT 87.345 99.405 92.690 99.840 ;
        RECT 92.865 99.405 94.075 100.495 ;
        RECT 94.245 99.405 94.535 100.570 ;
        RECT 98.110 99.840 98.460 101.090 ;
        RECT 103.630 99.840 103.980 101.090 ;
        RECT 106.435 100.495 106.955 101.035 ;
        RECT 94.705 99.405 100.050 99.840 ;
        RECT 100.225 99.405 105.570 99.840 ;
        RECT 105.745 99.405 106.955 100.495 ;
        RECT 107.125 99.405 107.415 100.570 ;
        RECT 110.990 99.840 111.340 101.090 ;
        RECT 116.510 99.840 116.860 101.090 ;
        RECT 119.315 100.495 119.835 101.035 ;
        RECT 107.585 99.405 112.930 99.840 ;
        RECT 113.105 99.405 118.450 99.840 ;
        RECT 118.625 99.405 119.835 100.495 ;
        RECT 120.005 99.405 120.295 100.570 ;
        RECT 123.870 99.840 124.220 101.090 ;
        RECT 129.390 99.840 129.740 101.090 ;
        RECT 132.195 100.495 132.715 101.035 ;
        RECT 120.465 99.405 125.810 99.840 ;
        RECT 125.985 99.405 131.330 99.840 ;
        RECT 131.505 99.405 132.715 100.495 ;
        RECT 132.885 99.405 133.175 100.570 ;
        RECT 136.750 99.840 137.100 101.090 ;
        RECT 140.685 100.495 142.375 101.015 ;
        RECT 133.345 99.405 138.690 99.840 ;
        RECT 138.865 99.405 142.375 100.495 ;
        RECT 143.005 100.495 143.525 101.035 ;
        RECT 143.005 99.405 144.215 100.495 ;
        RECT 55.520 99.235 144.300 99.405 ;
        RECT 55.605 98.145 56.815 99.235 ;
        RECT 56.985 98.800 62.330 99.235 ;
        RECT 62.505 98.800 67.850 99.235 ;
        RECT 56.295 97.605 56.815 98.145 ;
        RECT 60.390 97.550 60.740 98.800 ;
        RECT 65.910 97.550 66.260 98.800 ;
        RECT 68.485 98.070 68.775 99.235 ;
        RECT 68.945 98.800 74.290 99.235 ;
        RECT 74.465 98.800 79.810 99.235 ;
        RECT 79.985 98.800 85.330 99.235 ;
        RECT 85.505 98.800 90.850 99.235 ;
        RECT 72.350 97.550 72.700 98.800 ;
        RECT 77.870 97.550 78.220 98.800 ;
        RECT 83.390 97.550 83.740 98.800 ;
        RECT 88.910 97.550 89.260 98.800 ;
        RECT 91.025 98.145 93.615 99.235 ;
        RECT 92.405 97.625 93.615 98.145 ;
        RECT 94.245 98.070 94.535 99.235 ;
        RECT 94.705 98.800 100.050 99.235 ;
        RECT 100.225 98.800 105.570 99.235 ;
        RECT 105.745 98.800 111.090 99.235 ;
        RECT 111.265 98.800 116.610 99.235 ;
        RECT 98.110 97.550 98.460 98.800 ;
        RECT 103.630 97.550 103.980 98.800 ;
        RECT 109.150 97.550 109.500 98.800 ;
        RECT 114.670 97.550 115.020 98.800 ;
        RECT 116.785 98.145 119.375 99.235 ;
        RECT 118.165 97.625 119.375 98.145 ;
        RECT 120.005 98.070 120.295 99.235 ;
        RECT 120.465 98.800 125.810 99.235 ;
        RECT 125.985 98.800 131.330 99.235 ;
        RECT 131.505 98.800 136.850 99.235 ;
        RECT 137.025 98.800 142.370 99.235 ;
        RECT 123.870 97.550 124.220 98.800 ;
        RECT 129.390 97.550 129.740 98.800 ;
        RECT 134.910 97.550 135.260 98.800 ;
        RECT 140.430 97.550 140.780 98.800 ;
        RECT 143.005 98.145 144.215 99.235 ;
        RECT 143.005 97.605 143.525 98.145 ;
        RECT 56.295 95.055 56.815 95.595 ;
        RECT 55.605 93.965 56.815 95.055 ;
        RECT 60.390 94.400 60.740 95.650 ;
        RECT 65.910 94.400 66.260 95.650 ;
        RECT 71.430 94.400 71.780 95.650 ;
        RECT 76.950 94.400 77.300 95.650 ;
        RECT 79.985 95.055 80.735 95.575 ;
        RECT 56.985 93.965 62.330 94.400 ;
        RECT 62.505 93.965 67.850 94.400 ;
        RECT 68.025 93.965 73.370 94.400 ;
        RECT 73.545 93.965 78.890 94.400 ;
        RECT 79.065 93.965 80.735 95.055 ;
        RECT 81.365 93.965 81.655 95.130 ;
        RECT 85.230 94.400 85.580 95.650 ;
        RECT 90.750 94.400 91.100 95.650 ;
        RECT 96.270 94.400 96.620 95.650 ;
        RECT 101.790 94.400 102.140 95.650 ;
        RECT 105.285 95.055 106.495 95.575 ;
        RECT 81.825 93.965 87.170 94.400 ;
        RECT 87.345 93.965 92.690 94.400 ;
        RECT 92.865 93.965 98.210 94.400 ;
        RECT 98.385 93.965 103.730 94.400 ;
        RECT 103.905 93.965 106.495 95.055 ;
        RECT 107.125 93.965 107.415 95.130 ;
        RECT 110.990 94.400 111.340 95.650 ;
        RECT 116.510 94.400 116.860 95.650 ;
        RECT 122.030 94.400 122.380 95.650 ;
        RECT 127.550 94.400 127.900 95.650 ;
        RECT 131.045 95.055 132.255 95.575 ;
        RECT 107.585 93.965 112.930 94.400 ;
        RECT 113.105 93.965 118.450 94.400 ;
        RECT 118.625 93.965 123.970 94.400 ;
        RECT 124.145 93.965 129.490 94.400 ;
        RECT 129.665 93.965 132.255 95.055 ;
        RECT 132.885 93.965 133.175 95.130 ;
        RECT 136.750 94.400 137.100 95.650 ;
        RECT 140.685 95.055 142.375 95.575 ;
        RECT 133.345 93.965 138.690 94.400 ;
        RECT 138.865 93.965 142.375 95.055 ;
        RECT 143.005 95.055 143.525 95.595 ;
        RECT 143.005 93.965 144.215 95.055 ;
        RECT 55.520 93.795 144.300 93.965 ;
        RECT 55.605 92.705 56.815 93.795 ;
        RECT 56.985 93.360 62.330 93.795 ;
        RECT 62.505 93.360 67.850 93.795 ;
        RECT 56.295 92.165 56.815 92.705 ;
        RECT 60.390 92.110 60.740 93.360 ;
        RECT 65.910 92.110 66.260 93.360 ;
        RECT 68.485 92.630 68.775 93.795 ;
        RECT 68.945 93.360 74.290 93.795 ;
        RECT 74.465 93.360 79.810 93.795 ;
        RECT 79.985 93.360 85.330 93.795 ;
        RECT 85.505 93.360 90.850 93.795 ;
        RECT 72.350 92.110 72.700 93.360 ;
        RECT 77.870 92.110 78.220 93.360 ;
        RECT 83.390 92.110 83.740 93.360 ;
        RECT 88.910 92.110 89.260 93.360 ;
        RECT 91.025 92.705 93.615 93.795 ;
        RECT 92.405 92.185 93.615 92.705 ;
        RECT 94.245 92.630 94.535 93.795 ;
        RECT 94.705 93.360 100.050 93.795 ;
        RECT 100.225 93.360 105.570 93.795 ;
        RECT 105.745 93.360 111.090 93.795 ;
        RECT 111.265 93.360 116.610 93.795 ;
        RECT 98.110 92.110 98.460 93.360 ;
        RECT 103.630 92.110 103.980 93.360 ;
        RECT 109.150 92.110 109.500 93.360 ;
        RECT 114.670 92.110 115.020 93.360 ;
        RECT 116.785 92.705 119.375 93.795 ;
        RECT 118.165 92.185 119.375 92.705 ;
        RECT 120.005 92.630 120.295 93.795 ;
        RECT 120.465 93.360 125.810 93.795 ;
        RECT 125.985 93.360 131.330 93.795 ;
        RECT 131.505 93.360 136.850 93.795 ;
        RECT 137.025 93.360 142.370 93.795 ;
        RECT 123.870 92.110 124.220 93.360 ;
        RECT 129.390 92.110 129.740 93.360 ;
        RECT 134.910 92.110 135.260 93.360 ;
        RECT 140.430 92.110 140.780 93.360 ;
        RECT 143.005 92.705 144.215 93.795 ;
        RECT 143.005 92.165 143.525 92.705 ;
        RECT 56.295 89.615 56.815 90.155 ;
        RECT 55.605 88.525 56.815 89.615 ;
        RECT 60.390 88.960 60.740 90.210 ;
        RECT 65.910 88.960 66.260 90.210 ;
        RECT 71.430 88.960 71.780 90.210 ;
        RECT 76.950 88.960 77.300 90.210 ;
        RECT 79.985 89.615 80.735 90.135 ;
        RECT 56.985 88.525 62.330 88.960 ;
        RECT 62.505 88.525 67.850 88.960 ;
        RECT 68.025 88.525 73.370 88.960 ;
        RECT 73.545 88.525 78.890 88.960 ;
        RECT 79.065 88.525 80.735 89.615 ;
        RECT 81.365 88.525 81.655 89.690 ;
        RECT 85.230 88.960 85.580 90.210 ;
        RECT 90.750 88.960 91.100 90.210 ;
        RECT 96.270 88.960 96.620 90.210 ;
        RECT 101.790 88.960 102.140 90.210 ;
        RECT 105.285 89.615 106.495 90.135 ;
        RECT 81.825 88.525 87.170 88.960 ;
        RECT 87.345 88.525 92.690 88.960 ;
        RECT 92.865 88.525 98.210 88.960 ;
        RECT 98.385 88.525 103.730 88.960 ;
        RECT 103.905 88.525 106.495 89.615 ;
        RECT 107.125 88.525 107.415 89.690 ;
        RECT 110.990 88.960 111.340 90.210 ;
        RECT 116.510 88.960 116.860 90.210 ;
        RECT 122.030 88.960 122.380 90.210 ;
        RECT 127.550 88.960 127.900 90.210 ;
        RECT 131.045 89.615 132.255 90.135 ;
        RECT 107.585 88.525 112.930 88.960 ;
        RECT 113.105 88.525 118.450 88.960 ;
        RECT 118.625 88.525 123.970 88.960 ;
        RECT 124.145 88.525 129.490 88.960 ;
        RECT 129.665 88.525 132.255 89.615 ;
        RECT 132.885 88.525 133.175 89.690 ;
        RECT 136.750 88.960 137.100 90.210 ;
        RECT 140.685 89.615 142.375 90.135 ;
        RECT 133.345 88.525 138.690 88.960 ;
        RECT 138.865 88.525 142.375 89.615 ;
        RECT 143.005 89.615 143.525 90.155 ;
        RECT 143.005 88.525 144.215 89.615 ;
        RECT 55.520 88.355 144.300 88.525 ;
        RECT 55.605 87.265 56.815 88.355 ;
        RECT 56.985 87.920 62.330 88.355 ;
        RECT 62.505 87.920 67.850 88.355 ;
        RECT 56.295 86.725 56.815 87.265 ;
        RECT 60.390 86.670 60.740 87.920 ;
        RECT 65.910 86.670 66.260 87.920 ;
        RECT 68.485 87.190 68.775 88.355 ;
        RECT 68.945 87.920 74.290 88.355 ;
        RECT 74.465 87.920 79.810 88.355 ;
        RECT 79.985 87.920 85.330 88.355 ;
        RECT 85.505 87.920 90.850 88.355 ;
        RECT 72.350 86.670 72.700 87.920 ;
        RECT 77.870 86.670 78.220 87.920 ;
        RECT 83.390 86.670 83.740 87.920 ;
        RECT 88.910 86.670 89.260 87.920 ;
        RECT 91.025 87.265 93.615 88.355 ;
        RECT 92.405 86.745 93.615 87.265 ;
        RECT 94.245 87.190 94.535 88.355 ;
        RECT 94.705 87.920 100.050 88.355 ;
        RECT 100.225 87.920 105.570 88.355 ;
        RECT 105.745 87.920 111.090 88.355 ;
        RECT 111.265 87.920 116.610 88.355 ;
        RECT 98.110 86.670 98.460 87.920 ;
        RECT 103.630 86.670 103.980 87.920 ;
        RECT 109.150 86.670 109.500 87.920 ;
        RECT 114.670 86.670 115.020 87.920 ;
        RECT 116.785 87.265 119.375 88.355 ;
        RECT 118.165 86.745 119.375 87.265 ;
        RECT 120.005 87.190 120.295 88.355 ;
        RECT 120.465 87.920 125.810 88.355 ;
        RECT 125.985 87.920 131.330 88.355 ;
        RECT 131.505 87.920 136.850 88.355 ;
        RECT 137.025 87.920 142.370 88.355 ;
        RECT 123.870 86.670 124.220 87.920 ;
        RECT 129.390 86.670 129.740 87.920 ;
        RECT 134.910 86.670 135.260 87.920 ;
        RECT 140.430 86.670 140.780 87.920 ;
        RECT 143.005 87.265 144.215 88.355 ;
        RECT 143.005 86.725 143.525 87.265 ;
        RECT 56.295 84.175 56.815 84.715 ;
        RECT 55.605 83.085 56.815 84.175 ;
        RECT 60.390 83.520 60.740 84.770 ;
        RECT 65.910 83.520 66.260 84.770 ;
        RECT 71.430 83.520 71.780 84.770 ;
        RECT 76.950 83.520 77.300 84.770 ;
        RECT 79.985 84.175 80.735 84.695 ;
        RECT 56.985 83.085 62.330 83.520 ;
        RECT 62.505 83.085 67.850 83.520 ;
        RECT 68.025 83.085 73.370 83.520 ;
        RECT 73.545 83.085 78.890 83.520 ;
        RECT 79.065 83.085 80.735 84.175 ;
        RECT 81.365 83.085 81.655 84.250 ;
        RECT 85.230 83.520 85.580 84.770 ;
        RECT 90.750 83.520 91.100 84.770 ;
        RECT 96.270 83.520 96.620 84.770 ;
        RECT 101.790 83.520 102.140 84.770 ;
        RECT 105.285 84.175 106.495 84.695 ;
        RECT 81.825 83.085 87.170 83.520 ;
        RECT 87.345 83.085 92.690 83.520 ;
        RECT 92.865 83.085 98.210 83.520 ;
        RECT 98.385 83.085 103.730 83.520 ;
        RECT 103.905 83.085 106.495 84.175 ;
        RECT 107.125 83.085 107.415 84.250 ;
        RECT 110.990 83.520 111.340 84.770 ;
        RECT 116.510 83.520 116.860 84.770 ;
        RECT 122.030 83.520 122.380 84.770 ;
        RECT 127.550 83.520 127.900 84.770 ;
        RECT 131.045 84.175 132.255 84.695 ;
        RECT 107.585 83.085 112.930 83.520 ;
        RECT 113.105 83.085 118.450 83.520 ;
        RECT 118.625 83.085 123.970 83.520 ;
        RECT 124.145 83.085 129.490 83.520 ;
        RECT 129.665 83.085 132.255 84.175 ;
        RECT 132.885 83.085 133.175 84.250 ;
        RECT 136.750 83.520 137.100 84.770 ;
        RECT 140.685 84.175 142.375 84.695 ;
        RECT 133.345 83.085 138.690 83.520 ;
        RECT 138.865 83.085 142.375 84.175 ;
        RECT 143.005 84.175 143.525 84.715 ;
        RECT 143.005 83.085 144.215 84.175 ;
        RECT 55.520 82.915 144.300 83.085 ;
        RECT 55.605 81.825 56.815 82.915 ;
        RECT 56.985 82.480 62.330 82.915 ;
        RECT 62.505 82.480 67.850 82.915 ;
        RECT 56.295 81.285 56.815 81.825 ;
        RECT 60.390 81.230 60.740 82.480 ;
        RECT 65.910 81.230 66.260 82.480 ;
        RECT 68.485 81.750 68.775 82.915 ;
        RECT 68.945 82.480 74.290 82.915 ;
        RECT 74.465 82.480 79.810 82.915 ;
        RECT 79.985 82.480 85.330 82.915 ;
        RECT 85.505 82.480 90.850 82.915 ;
        RECT 72.350 81.230 72.700 82.480 ;
        RECT 77.870 81.230 78.220 82.480 ;
        RECT 83.390 81.230 83.740 82.480 ;
        RECT 88.910 81.230 89.260 82.480 ;
        RECT 91.025 81.825 93.615 82.915 ;
        RECT 92.405 81.305 93.615 81.825 ;
        RECT 94.245 81.750 94.535 82.915 ;
        RECT 94.705 82.480 100.050 82.915 ;
        RECT 100.225 82.480 105.570 82.915 ;
        RECT 105.745 82.480 111.090 82.915 ;
        RECT 111.265 82.480 116.610 82.915 ;
        RECT 98.110 81.230 98.460 82.480 ;
        RECT 103.630 81.230 103.980 82.480 ;
        RECT 109.150 81.230 109.500 82.480 ;
        RECT 114.670 81.230 115.020 82.480 ;
        RECT 116.785 81.825 119.375 82.915 ;
        RECT 118.165 81.305 119.375 81.825 ;
        RECT 120.005 81.750 120.295 82.915 ;
        RECT 120.465 82.480 125.810 82.915 ;
        RECT 125.985 82.480 131.330 82.915 ;
        RECT 131.505 82.480 136.850 82.915 ;
        RECT 137.025 82.480 142.370 82.915 ;
        RECT 123.870 81.230 124.220 82.480 ;
        RECT 129.390 81.230 129.740 82.480 ;
        RECT 134.910 81.230 135.260 82.480 ;
        RECT 140.430 81.230 140.780 82.480 ;
        RECT 143.005 81.825 144.215 82.915 ;
        RECT 143.005 81.285 143.525 81.825 ;
        RECT 56.295 78.735 56.815 79.275 ;
        RECT 55.605 77.645 56.815 78.735 ;
        RECT 60.390 78.080 60.740 79.330 ;
        RECT 65.910 78.080 66.260 79.330 ;
        RECT 71.430 78.080 71.780 79.330 ;
        RECT 76.950 78.080 77.300 79.330 ;
        RECT 79.985 78.735 80.735 79.255 ;
        RECT 56.985 77.645 62.330 78.080 ;
        RECT 62.505 77.645 67.850 78.080 ;
        RECT 68.025 77.645 73.370 78.080 ;
        RECT 73.545 77.645 78.890 78.080 ;
        RECT 79.065 77.645 80.735 78.735 ;
        RECT 81.365 77.645 81.655 78.810 ;
        RECT 85.230 78.080 85.580 79.330 ;
        RECT 90.750 78.080 91.100 79.330 ;
        RECT 96.270 78.080 96.620 79.330 ;
        RECT 101.790 78.080 102.140 79.330 ;
        RECT 105.285 78.735 106.495 79.255 ;
        RECT 81.825 77.645 87.170 78.080 ;
        RECT 87.345 77.645 92.690 78.080 ;
        RECT 92.865 77.645 98.210 78.080 ;
        RECT 98.385 77.645 103.730 78.080 ;
        RECT 103.905 77.645 106.495 78.735 ;
        RECT 107.125 77.645 107.415 78.810 ;
        RECT 110.990 78.080 111.340 79.330 ;
        RECT 116.510 78.080 116.860 79.330 ;
        RECT 122.030 78.080 122.380 79.330 ;
        RECT 127.550 78.080 127.900 79.330 ;
        RECT 131.045 78.735 132.255 79.255 ;
        RECT 107.585 77.645 112.930 78.080 ;
        RECT 113.105 77.645 118.450 78.080 ;
        RECT 118.625 77.645 123.970 78.080 ;
        RECT 124.145 77.645 129.490 78.080 ;
        RECT 129.665 77.645 132.255 78.735 ;
        RECT 132.885 77.645 133.175 78.810 ;
        RECT 136.750 78.080 137.100 79.330 ;
        RECT 140.685 78.735 142.375 79.255 ;
        RECT 133.345 77.645 138.690 78.080 ;
        RECT 138.865 77.645 142.375 78.735 ;
        RECT 143.005 78.735 143.525 79.275 ;
        RECT 143.005 77.645 144.215 78.735 ;
        RECT 55.520 77.475 144.300 77.645 ;
        RECT 55.605 76.385 56.815 77.475 ;
        RECT 56.985 77.040 62.330 77.475 ;
        RECT 62.505 77.040 67.850 77.475 ;
        RECT 56.295 75.845 56.815 76.385 ;
        RECT 60.390 75.790 60.740 77.040 ;
        RECT 65.910 75.790 66.260 77.040 ;
        RECT 68.485 76.310 68.775 77.475 ;
        RECT 68.945 77.040 74.290 77.475 ;
        RECT 74.465 77.040 79.810 77.475 ;
        RECT 79.985 77.040 85.330 77.475 ;
        RECT 85.505 77.040 90.850 77.475 ;
        RECT 72.350 75.790 72.700 77.040 ;
        RECT 77.870 75.790 78.220 77.040 ;
        RECT 83.390 75.790 83.740 77.040 ;
        RECT 88.910 75.790 89.260 77.040 ;
        RECT 91.025 76.385 93.615 77.475 ;
        RECT 92.405 75.865 93.615 76.385 ;
        RECT 94.245 76.310 94.535 77.475 ;
        RECT 94.705 77.040 100.050 77.475 ;
        RECT 100.225 77.040 105.570 77.475 ;
        RECT 105.745 77.040 111.090 77.475 ;
        RECT 111.265 77.040 116.610 77.475 ;
        RECT 98.110 75.790 98.460 77.040 ;
        RECT 103.630 75.790 103.980 77.040 ;
        RECT 109.150 75.790 109.500 77.040 ;
        RECT 114.670 75.790 115.020 77.040 ;
        RECT 116.785 76.385 119.375 77.475 ;
        RECT 118.165 75.865 119.375 76.385 ;
        RECT 120.005 76.310 120.295 77.475 ;
        RECT 120.465 77.040 125.810 77.475 ;
        RECT 125.985 77.040 131.330 77.475 ;
        RECT 131.505 77.040 136.850 77.475 ;
        RECT 137.025 77.040 142.370 77.475 ;
        RECT 123.870 75.790 124.220 77.040 ;
        RECT 129.390 75.790 129.740 77.040 ;
        RECT 134.910 75.790 135.260 77.040 ;
        RECT 140.430 75.790 140.780 77.040 ;
        RECT 143.005 76.385 144.215 77.475 ;
        RECT 143.005 75.845 143.525 76.385 ;
        RECT 56.295 73.295 56.815 73.835 ;
        RECT 55.605 72.205 56.815 73.295 ;
        RECT 60.390 72.640 60.740 73.890 ;
        RECT 65.910 72.640 66.260 73.890 ;
        RECT 68.945 73.295 69.695 73.815 ;
        RECT 56.985 72.205 62.330 72.640 ;
        RECT 62.505 72.205 67.850 72.640 ;
        RECT 68.025 72.205 69.695 73.295 ;
        RECT 70.365 72.205 70.595 73.345 ;
        RECT 71.265 72.205 71.475 73.345 ;
        RECT 72.180 72.205 72.510 72.965 ;
        RECT 73.110 72.205 73.370 73.355 ;
        RECT 76.950 72.640 77.300 73.890 ;
        RECT 79.985 73.295 80.735 73.815 ;
        RECT 73.545 72.205 78.890 72.640 ;
        RECT 79.065 72.205 80.735 73.295 ;
        RECT 81.365 72.205 81.655 73.370 ;
        RECT 85.230 72.640 85.580 73.890 ;
        RECT 90.750 72.640 91.100 73.890 ;
        RECT 96.270 72.640 96.620 73.890 ;
        RECT 101.790 72.640 102.140 73.890 ;
        RECT 105.285 73.295 106.495 73.815 ;
        RECT 81.825 72.205 87.170 72.640 ;
        RECT 87.345 72.205 92.690 72.640 ;
        RECT 92.865 72.205 98.210 72.640 ;
        RECT 98.385 72.205 103.730 72.640 ;
        RECT 103.905 72.205 106.495 73.295 ;
        RECT 107.125 72.205 107.415 73.370 ;
        RECT 110.990 72.640 111.340 73.890 ;
        RECT 116.510 72.640 116.860 73.890 ;
        RECT 122.030 72.640 122.380 73.890 ;
        RECT 127.550 72.640 127.900 73.890 ;
        RECT 131.045 73.295 132.255 73.815 ;
        RECT 107.585 72.205 112.930 72.640 ;
        RECT 113.105 72.205 118.450 72.640 ;
        RECT 118.625 72.205 123.970 72.640 ;
        RECT 124.145 72.205 129.490 72.640 ;
        RECT 129.665 72.205 132.255 73.295 ;
        RECT 132.885 72.205 133.175 73.370 ;
        RECT 136.750 72.640 137.100 73.890 ;
        RECT 140.685 73.295 142.375 73.815 ;
        RECT 133.345 72.205 138.690 72.640 ;
        RECT 138.865 72.205 142.375 73.295 ;
        RECT 143.005 73.295 143.525 73.835 ;
        RECT 143.005 72.205 144.215 73.295 ;
        RECT 55.520 72.035 144.300 72.205 ;
        RECT 55.605 70.945 56.815 72.035 ;
        RECT 56.985 70.945 60.495 72.035 ;
        RECT 56.295 70.405 56.815 70.945 ;
        RECT 58.805 70.425 60.495 70.945 ;
        RECT 61.185 70.895 61.395 72.035 ;
        RECT 62.065 70.895 62.295 72.035 ;
        RECT 62.505 70.895 62.785 72.035 ;
        RECT 63.455 70.895 63.715 72.035 ;
        RECT 65.675 71.575 66.040 72.035 ;
        RECT 66.635 71.575 66.965 72.035 ;
        RECT 68.485 70.870 68.775 72.035 ;
        RECT 68.945 71.600 74.290 72.035 ;
        RECT 74.465 71.600 79.810 72.035 ;
        RECT 79.985 71.600 85.330 72.035 ;
        RECT 85.505 71.600 90.850 72.035 ;
        RECT 72.350 70.350 72.700 71.600 ;
        RECT 77.870 70.350 78.220 71.600 ;
        RECT 83.390 70.350 83.740 71.600 ;
        RECT 88.910 70.350 89.260 71.600 ;
        RECT 91.025 70.945 93.615 72.035 ;
        RECT 92.405 70.425 93.615 70.945 ;
        RECT 94.245 70.870 94.535 72.035 ;
        RECT 94.705 71.600 100.050 72.035 ;
        RECT 100.225 71.600 105.570 72.035 ;
        RECT 105.745 71.600 111.090 72.035 ;
        RECT 111.265 71.600 116.610 72.035 ;
        RECT 98.110 70.350 98.460 71.600 ;
        RECT 103.630 70.350 103.980 71.600 ;
        RECT 109.150 70.350 109.500 71.600 ;
        RECT 114.670 70.350 115.020 71.600 ;
        RECT 116.785 70.945 119.375 72.035 ;
        RECT 118.165 70.425 119.375 70.945 ;
        RECT 120.005 70.870 120.295 72.035 ;
        RECT 120.465 71.600 125.810 72.035 ;
        RECT 125.985 71.600 131.330 72.035 ;
        RECT 131.505 71.600 136.850 72.035 ;
        RECT 137.025 71.600 142.370 72.035 ;
        RECT 123.870 70.350 124.220 71.600 ;
        RECT 129.390 70.350 129.740 71.600 ;
        RECT 134.910 70.350 135.260 71.600 ;
        RECT 140.430 70.350 140.780 71.600 ;
        RECT 143.005 70.945 144.215 72.035 ;
        RECT 143.005 70.405 143.525 70.945 ;
        RECT 56.295 67.855 56.815 68.395 ;
        RECT 55.605 66.765 56.815 67.855 ;
        RECT 57.425 66.765 57.755 67.525 ;
        RECT 61.770 67.200 62.120 68.450 ;
        RECT 58.365 66.765 63.710 67.200 ;
        RECT 64.805 66.765 65.065 67.905 ;
        RECT 65.735 66.765 65.905 67.565 ;
        RECT 66.575 66.765 66.830 67.565 ;
        RECT 67.535 66.765 67.970 67.555 ;
        RECT 74.650 67.200 75.000 68.450 ;
        RECT 78.585 67.855 80.275 68.375 ;
        RECT 69.000 66.765 69.330 67.125 ;
        RECT 71.245 66.765 76.590 67.200 ;
        RECT 76.765 66.765 80.275 67.855 ;
        RECT 81.365 66.765 81.655 67.930 ;
        RECT 85.230 67.200 85.580 68.450 ;
        RECT 90.750 67.200 91.100 68.450 ;
        RECT 96.270 67.200 96.620 68.450 ;
        RECT 101.790 67.200 102.140 68.450 ;
        RECT 105.285 67.855 106.495 68.375 ;
        RECT 81.825 66.765 87.170 67.200 ;
        RECT 87.345 66.765 92.690 67.200 ;
        RECT 92.865 66.765 98.210 67.200 ;
        RECT 98.385 66.765 103.730 67.200 ;
        RECT 103.905 66.765 106.495 67.855 ;
        RECT 107.125 66.765 107.415 67.930 ;
        RECT 110.990 67.200 111.340 68.450 ;
        RECT 116.510 67.200 116.860 68.450 ;
        RECT 122.030 67.200 122.380 68.450 ;
        RECT 127.550 67.200 127.900 68.450 ;
        RECT 131.045 67.855 132.255 68.375 ;
        RECT 107.585 66.765 112.930 67.200 ;
        RECT 113.105 66.765 118.450 67.200 ;
        RECT 118.625 66.765 123.970 67.200 ;
        RECT 124.145 66.765 129.490 67.200 ;
        RECT 129.665 66.765 132.255 67.855 ;
        RECT 132.885 66.765 133.175 67.930 ;
        RECT 136.750 67.200 137.100 68.450 ;
        RECT 140.685 67.855 142.375 68.375 ;
        RECT 133.345 66.765 138.690 67.200 ;
        RECT 138.865 66.765 142.375 67.855 ;
        RECT 143.005 67.855 143.525 68.395 ;
        RECT 143.005 66.765 144.215 67.855 ;
        RECT 55.520 66.595 144.300 66.765 ;
        RECT 55.605 65.505 56.815 66.595 ;
        RECT 57.425 65.835 57.755 66.595 ;
        RECT 58.365 66.160 63.710 66.595 ;
        RECT 56.295 64.965 56.815 65.505 ;
        RECT 61.770 64.910 62.120 66.160 ;
        RECT 63.885 65.505 67.395 66.595 ;
        RECT 65.705 64.985 67.395 65.505 ;
        RECT 68.485 65.430 68.775 66.595 ;
        RECT 68.945 66.160 74.290 66.595 ;
        RECT 74.465 66.160 79.810 66.595 ;
        RECT 79.985 66.160 85.330 66.595 ;
        RECT 85.505 66.160 90.850 66.595 ;
        RECT 72.350 64.910 72.700 66.160 ;
        RECT 77.870 64.910 78.220 66.160 ;
        RECT 83.390 64.910 83.740 66.160 ;
        RECT 88.910 64.910 89.260 66.160 ;
        RECT 91.025 65.505 93.615 66.595 ;
        RECT 92.405 64.985 93.615 65.505 ;
        RECT 94.245 65.430 94.535 66.595 ;
        RECT 94.705 66.160 100.050 66.595 ;
        RECT 100.225 66.160 105.570 66.595 ;
        RECT 105.745 66.160 111.090 66.595 ;
        RECT 111.265 66.160 116.610 66.595 ;
        RECT 98.110 64.910 98.460 66.160 ;
        RECT 103.630 64.910 103.980 66.160 ;
        RECT 109.150 64.910 109.500 66.160 ;
        RECT 114.670 64.910 115.020 66.160 ;
        RECT 116.785 65.505 119.375 66.595 ;
        RECT 118.165 64.985 119.375 65.505 ;
        RECT 120.005 65.430 120.295 66.595 ;
        RECT 120.465 66.160 125.810 66.595 ;
        RECT 125.985 66.160 131.330 66.595 ;
        RECT 131.505 66.160 136.850 66.595 ;
        RECT 137.025 66.160 142.370 66.595 ;
        RECT 123.870 64.910 124.220 66.160 ;
        RECT 129.390 64.910 129.740 66.160 ;
        RECT 134.910 64.910 135.260 66.160 ;
        RECT 140.430 64.910 140.780 66.160 ;
        RECT 143.005 65.505 144.215 66.595 ;
        RECT 143.005 64.965 143.525 65.505 ;
        RECT 56.295 62.415 56.815 62.955 ;
        RECT 55.605 61.325 56.815 62.415 ;
        RECT 60.390 61.760 60.740 63.010 ;
        RECT 63.885 62.415 65.095 62.935 ;
        RECT 56.985 61.325 62.330 61.760 ;
        RECT 62.505 61.325 65.095 62.415 ;
        RECT 66.165 61.325 66.495 62.085 ;
        RECT 70.510 61.760 70.860 63.010 ;
        RECT 76.030 61.760 76.380 63.010 ;
        RECT 79.525 62.415 80.735 62.935 ;
        RECT 67.105 61.325 72.450 61.760 ;
        RECT 72.625 61.325 77.970 61.760 ;
        RECT 78.145 61.325 80.735 62.415 ;
        RECT 81.365 61.325 81.655 62.490 ;
        RECT 85.230 61.760 85.580 63.010 ;
        RECT 90.750 61.760 91.100 63.010 ;
        RECT 96.270 61.760 96.620 63.010 ;
        RECT 101.790 61.760 102.140 63.010 ;
        RECT 105.285 62.415 106.495 62.935 ;
        RECT 81.825 61.325 87.170 61.760 ;
        RECT 87.345 61.325 92.690 61.760 ;
        RECT 92.865 61.325 98.210 61.760 ;
        RECT 98.385 61.325 103.730 61.760 ;
        RECT 103.905 61.325 106.495 62.415 ;
        RECT 107.125 61.325 107.415 62.490 ;
        RECT 110.990 61.760 111.340 63.010 ;
        RECT 116.510 61.760 116.860 63.010 ;
        RECT 122.030 61.760 122.380 63.010 ;
        RECT 127.550 61.760 127.900 63.010 ;
        RECT 131.045 62.415 132.255 62.935 ;
        RECT 107.585 61.325 112.930 61.760 ;
        RECT 113.105 61.325 118.450 61.760 ;
        RECT 118.625 61.325 123.970 61.760 ;
        RECT 124.145 61.325 129.490 61.760 ;
        RECT 129.665 61.325 132.255 62.415 ;
        RECT 132.885 61.325 133.175 62.490 ;
        RECT 136.750 61.760 137.100 63.010 ;
        RECT 140.685 62.415 142.375 62.935 ;
        RECT 133.345 61.325 138.690 61.760 ;
        RECT 138.865 61.325 142.375 62.415 ;
        RECT 143.005 62.415 143.525 62.955 ;
        RECT 143.005 61.325 144.215 62.415 ;
        RECT 55.520 61.155 144.300 61.325 ;
        RECT 55.605 60.065 56.815 61.155 ;
        RECT 56.985 60.720 62.330 61.155 ;
        RECT 56.295 59.525 56.815 60.065 ;
        RECT 60.390 59.470 60.740 60.720 ;
        RECT 62.505 60.065 66.015 61.155 ;
        RECT 64.325 59.545 66.015 60.065 ;
        RECT 66.645 60.015 66.905 61.155 ;
        RECT 67.575 60.015 67.855 61.155 ;
        RECT 68.485 59.990 68.775 61.155 ;
        RECT 68.945 60.720 74.290 61.155 ;
        RECT 74.465 60.720 79.810 61.155 ;
        RECT 79.985 60.720 85.330 61.155 ;
        RECT 85.505 60.720 90.850 61.155 ;
        RECT 72.350 59.470 72.700 60.720 ;
        RECT 77.870 59.470 78.220 60.720 ;
        RECT 83.390 59.470 83.740 60.720 ;
        RECT 88.910 59.470 89.260 60.720 ;
        RECT 91.025 60.065 93.615 61.155 ;
        RECT 92.405 59.545 93.615 60.065 ;
        RECT 94.245 59.990 94.535 61.155 ;
        RECT 94.705 60.720 100.050 61.155 ;
        RECT 100.225 60.720 105.570 61.155 ;
        RECT 105.745 60.720 111.090 61.155 ;
        RECT 111.265 60.720 116.610 61.155 ;
        RECT 98.110 59.470 98.460 60.720 ;
        RECT 103.630 59.470 103.980 60.720 ;
        RECT 109.150 59.470 109.500 60.720 ;
        RECT 114.670 59.470 115.020 60.720 ;
        RECT 116.785 60.065 119.375 61.155 ;
        RECT 118.165 59.545 119.375 60.065 ;
        RECT 120.005 59.990 120.295 61.155 ;
        RECT 120.465 60.720 125.810 61.155 ;
        RECT 125.985 60.720 131.330 61.155 ;
        RECT 131.505 60.720 136.850 61.155 ;
        RECT 137.025 60.720 142.370 61.155 ;
        RECT 123.870 59.470 124.220 60.720 ;
        RECT 129.390 59.470 129.740 60.720 ;
        RECT 134.910 59.470 135.260 60.720 ;
        RECT 140.430 59.470 140.780 60.720 ;
        RECT 143.005 60.065 144.215 61.155 ;
        RECT 143.005 59.525 143.525 60.065 ;
        RECT 56.295 56.975 56.815 57.515 ;
        RECT 58.805 56.975 60.495 57.495 ;
        RECT 55.605 55.885 56.815 56.975 ;
        RECT 56.985 55.885 60.495 56.975 ;
        RECT 62.335 55.885 62.505 56.645 ;
        RECT 64.875 55.885 65.045 57.025 ;
        RECT 66.235 55.885 66.405 57.025 ;
        RECT 68.775 55.885 68.945 56.645 ;
        RECT 69.905 55.885 70.135 57.025 ;
        RECT 70.805 55.885 71.015 57.025 ;
        RECT 71.285 55.885 71.515 57.025 ;
        RECT 72.185 55.885 72.395 57.025 ;
        RECT 76.030 56.320 76.380 57.570 ;
        RECT 79.525 56.975 80.735 57.495 ;
        RECT 72.625 55.885 77.970 56.320 ;
        RECT 78.145 55.885 80.735 56.975 ;
        RECT 81.365 55.885 81.655 57.050 ;
        RECT 85.230 56.320 85.580 57.570 ;
        RECT 90.750 56.320 91.100 57.570 ;
        RECT 96.270 56.320 96.620 57.570 ;
        RECT 101.790 56.320 102.140 57.570 ;
        RECT 105.285 56.975 106.495 57.495 ;
        RECT 81.825 55.885 87.170 56.320 ;
        RECT 87.345 55.885 92.690 56.320 ;
        RECT 92.865 55.885 98.210 56.320 ;
        RECT 98.385 55.885 103.730 56.320 ;
        RECT 103.905 55.885 106.495 56.975 ;
        RECT 107.125 55.885 107.415 57.050 ;
        RECT 110.990 56.320 111.340 57.570 ;
        RECT 116.510 56.320 116.860 57.570 ;
        RECT 122.030 56.320 122.380 57.570 ;
        RECT 127.550 56.320 127.900 57.570 ;
        RECT 131.045 56.975 132.255 57.495 ;
        RECT 107.585 55.885 112.930 56.320 ;
        RECT 113.105 55.885 118.450 56.320 ;
        RECT 118.625 55.885 123.970 56.320 ;
        RECT 124.145 55.885 129.490 56.320 ;
        RECT 129.665 55.885 132.255 56.975 ;
        RECT 132.885 55.885 133.175 57.050 ;
        RECT 136.750 56.320 137.100 57.570 ;
        RECT 140.685 56.975 142.375 57.495 ;
        RECT 133.345 55.885 138.690 56.320 ;
        RECT 138.865 55.885 142.375 56.975 ;
        RECT 143.005 56.975 143.525 57.515 ;
        RECT 143.005 55.885 144.215 56.975 ;
        RECT 55.520 55.715 144.300 55.885 ;
        RECT 55.605 54.625 56.815 55.715 ;
        RECT 56.985 55.280 62.330 55.715 ;
        RECT 56.295 54.085 56.815 54.625 ;
        RECT 60.390 54.030 60.740 55.280 ;
        RECT 62.505 54.625 65.095 55.715 ;
        RECT 65.705 54.955 66.035 55.715 ;
        RECT 63.885 54.105 65.095 54.625 ;
        RECT 66.685 54.575 66.915 55.715 ;
        RECT 67.585 54.575 67.795 55.715 ;
        RECT 68.485 54.550 68.775 55.715 ;
        RECT 68.945 55.280 74.290 55.715 ;
        RECT 74.465 55.280 79.810 55.715 ;
        RECT 79.985 55.280 85.330 55.715 ;
        RECT 85.505 55.280 90.850 55.715 ;
        RECT 72.350 54.030 72.700 55.280 ;
        RECT 77.870 54.030 78.220 55.280 ;
        RECT 83.390 54.030 83.740 55.280 ;
        RECT 88.910 54.030 89.260 55.280 ;
        RECT 91.025 54.625 93.615 55.715 ;
        RECT 92.405 54.105 93.615 54.625 ;
        RECT 94.245 54.550 94.535 55.715 ;
        RECT 94.705 55.280 100.050 55.715 ;
        RECT 100.225 55.280 105.570 55.715 ;
        RECT 105.745 55.280 111.090 55.715 ;
        RECT 111.265 55.280 116.610 55.715 ;
        RECT 98.110 54.030 98.460 55.280 ;
        RECT 103.630 54.030 103.980 55.280 ;
        RECT 109.150 54.030 109.500 55.280 ;
        RECT 114.670 54.030 115.020 55.280 ;
        RECT 116.785 54.625 119.375 55.715 ;
        RECT 118.165 54.105 119.375 54.625 ;
        RECT 120.005 54.550 120.295 55.715 ;
        RECT 120.465 55.280 125.810 55.715 ;
        RECT 125.985 55.280 131.330 55.715 ;
        RECT 131.505 55.280 136.850 55.715 ;
        RECT 137.025 55.280 142.370 55.715 ;
        RECT 123.870 54.030 124.220 55.280 ;
        RECT 129.390 54.030 129.740 55.280 ;
        RECT 134.910 54.030 135.260 55.280 ;
        RECT 140.430 54.030 140.780 55.280 ;
        RECT 143.005 54.625 144.215 55.715 ;
        RECT 143.005 54.085 143.525 54.625 ;
        RECT 56.295 51.535 56.815 52.075 ;
        RECT 55.605 50.445 56.815 51.535 ;
        RECT 60.390 50.880 60.740 52.130 ;
        RECT 65.910 50.880 66.260 52.130 ;
        RECT 71.430 50.880 71.780 52.130 ;
        RECT 76.950 50.880 77.300 52.130 ;
        RECT 79.985 51.535 80.735 52.055 ;
        RECT 56.985 50.445 62.330 50.880 ;
        RECT 62.505 50.445 67.850 50.880 ;
        RECT 68.025 50.445 73.370 50.880 ;
        RECT 73.545 50.445 78.890 50.880 ;
        RECT 79.065 50.445 80.735 51.535 ;
        RECT 81.365 50.445 81.655 51.610 ;
        RECT 85.230 50.880 85.580 52.130 ;
        RECT 90.750 50.880 91.100 52.130 ;
        RECT 96.270 50.880 96.620 52.130 ;
        RECT 101.790 50.880 102.140 52.130 ;
        RECT 105.285 51.535 106.495 52.055 ;
        RECT 81.825 50.445 87.170 50.880 ;
        RECT 87.345 50.445 92.690 50.880 ;
        RECT 92.865 50.445 98.210 50.880 ;
        RECT 98.385 50.445 103.730 50.880 ;
        RECT 103.905 50.445 106.495 51.535 ;
        RECT 107.125 50.445 107.415 51.610 ;
        RECT 110.990 50.880 111.340 52.130 ;
        RECT 116.510 50.880 116.860 52.130 ;
        RECT 122.030 50.880 122.380 52.130 ;
        RECT 127.550 50.880 127.900 52.130 ;
        RECT 131.045 51.535 132.255 52.055 ;
        RECT 107.585 50.445 112.930 50.880 ;
        RECT 113.105 50.445 118.450 50.880 ;
        RECT 118.625 50.445 123.970 50.880 ;
        RECT 124.145 50.445 129.490 50.880 ;
        RECT 129.665 50.445 132.255 51.535 ;
        RECT 132.885 50.445 133.175 51.610 ;
        RECT 136.750 50.880 137.100 52.130 ;
        RECT 140.685 51.535 142.375 52.055 ;
        RECT 133.345 50.445 138.690 50.880 ;
        RECT 138.865 50.445 142.375 51.535 ;
        RECT 143.005 51.535 143.525 52.075 ;
        RECT 143.005 50.445 144.215 51.535 ;
        RECT 55.520 50.275 144.300 50.445 ;
        RECT 55.605 49.185 56.815 50.275 ;
        RECT 56.985 49.840 62.330 50.275 ;
        RECT 62.505 49.840 67.850 50.275 ;
        RECT 56.295 48.645 56.815 49.185 ;
        RECT 60.390 48.590 60.740 49.840 ;
        RECT 65.910 48.590 66.260 49.840 ;
        RECT 68.485 49.110 68.775 50.275 ;
        RECT 68.945 49.840 74.290 50.275 ;
        RECT 74.465 49.840 79.810 50.275 ;
        RECT 79.985 49.840 85.330 50.275 ;
        RECT 85.505 49.840 90.850 50.275 ;
        RECT 72.350 48.590 72.700 49.840 ;
        RECT 77.870 48.590 78.220 49.840 ;
        RECT 83.390 48.590 83.740 49.840 ;
        RECT 88.910 48.590 89.260 49.840 ;
        RECT 91.025 49.185 93.615 50.275 ;
        RECT 92.405 48.665 93.615 49.185 ;
        RECT 94.245 49.110 94.535 50.275 ;
        RECT 94.705 49.840 100.050 50.275 ;
        RECT 100.225 49.840 105.570 50.275 ;
        RECT 105.745 49.840 111.090 50.275 ;
        RECT 111.265 49.840 116.610 50.275 ;
        RECT 98.110 48.590 98.460 49.840 ;
        RECT 103.630 48.590 103.980 49.840 ;
        RECT 109.150 48.590 109.500 49.840 ;
        RECT 114.670 48.590 115.020 49.840 ;
        RECT 116.785 49.185 119.375 50.275 ;
        RECT 118.165 48.665 119.375 49.185 ;
        RECT 120.005 49.110 120.295 50.275 ;
        RECT 120.465 49.840 125.810 50.275 ;
        RECT 125.985 49.840 131.330 50.275 ;
        RECT 131.505 49.840 136.850 50.275 ;
        RECT 137.025 49.840 142.370 50.275 ;
        RECT 123.870 48.590 124.220 49.840 ;
        RECT 129.390 48.590 129.740 49.840 ;
        RECT 134.910 48.590 135.260 49.840 ;
        RECT 140.430 48.590 140.780 49.840 ;
        RECT 143.005 49.185 144.215 50.275 ;
        RECT 143.005 48.645 143.525 49.185 ;
        RECT 56.295 46.095 56.815 46.635 ;
        RECT 55.605 45.005 56.815 46.095 ;
        RECT 60.390 45.440 60.740 46.690 ;
        RECT 65.910 45.440 66.260 46.690 ;
        RECT 71.430 45.440 71.780 46.690 ;
        RECT 76.950 45.440 77.300 46.690 ;
        RECT 79.985 46.095 80.735 46.615 ;
        RECT 56.985 45.005 62.330 45.440 ;
        RECT 62.505 45.005 67.850 45.440 ;
        RECT 68.025 45.005 73.370 45.440 ;
        RECT 73.545 45.005 78.890 45.440 ;
        RECT 79.065 45.005 80.735 46.095 ;
        RECT 81.365 45.005 81.655 46.170 ;
        RECT 85.230 45.440 85.580 46.690 ;
        RECT 90.750 45.440 91.100 46.690 ;
        RECT 96.270 45.440 96.620 46.690 ;
        RECT 101.790 45.440 102.140 46.690 ;
        RECT 105.285 46.095 106.495 46.615 ;
        RECT 81.825 45.005 87.170 45.440 ;
        RECT 87.345 45.005 92.690 45.440 ;
        RECT 92.865 45.005 98.210 45.440 ;
        RECT 98.385 45.005 103.730 45.440 ;
        RECT 103.905 45.005 106.495 46.095 ;
        RECT 107.125 45.005 107.415 46.170 ;
        RECT 110.990 45.440 111.340 46.690 ;
        RECT 116.510 45.440 116.860 46.690 ;
        RECT 122.030 45.440 122.380 46.690 ;
        RECT 127.550 45.440 127.900 46.690 ;
        RECT 131.045 46.095 132.255 46.615 ;
        RECT 107.585 45.005 112.930 45.440 ;
        RECT 113.105 45.005 118.450 45.440 ;
        RECT 118.625 45.005 123.970 45.440 ;
        RECT 124.145 45.005 129.490 45.440 ;
        RECT 129.665 45.005 132.255 46.095 ;
        RECT 132.885 45.005 133.175 46.170 ;
        RECT 136.750 45.440 137.100 46.690 ;
        RECT 140.685 46.095 142.375 46.615 ;
        RECT 133.345 45.005 138.690 45.440 ;
        RECT 138.865 45.005 142.375 46.095 ;
        RECT 143.005 46.095 143.525 46.635 ;
        RECT 143.005 45.005 144.215 46.095 ;
        RECT 55.520 44.835 144.300 45.005 ;
        RECT 55.605 43.745 56.815 44.835 ;
        RECT 56.985 44.400 62.330 44.835 ;
        RECT 62.505 44.400 67.850 44.835 ;
        RECT 56.295 43.205 56.815 43.745 ;
        RECT 60.390 43.150 60.740 44.400 ;
        RECT 65.910 43.150 66.260 44.400 ;
        RECT 68.485 43.670 68.775 44.835 ;
        RECT 68.945 44.400 74.290 44.835 ;
        RECT 74.465 44.400 79.810 44.835 ;
        RECT 79.985 44.400 85.330 44.835 ;
        RECT 85.505 44.400 90.850 44.835 ;
        RECT 72.350 43.150 72.700 44.400 ;
        RECT 77.870 43.150 78.220 44.400 ;
        RECT 83.390 43.150 83.740 44.400 ;
        RECT 88.910 43.150 89.260 44.400 ;
        RECT 91.025 43.745 93.615 44.835 ;
        RECT 92.405 43.225 93.615 43.745 ;
        RECT 94.245 43.670 94.535 44.835 ;
        RECT 94.705 44.400 100.050 44.835 ;
        RECT 100.225 44.400 105.570 44.835 ;
        RECT 105.745 44.400 111.090 44.835 ;
        RECT 111.265 44.400 116.610 44.835 ;
        RECT 98.110 43.150 98.460 44.400 ;
        RECT 103.630 43.150 103.980 44.400 ;
        RECT 109.150 43.150 109.500 44.400 ;
        RECT 114.670 43.150 115.020 44.400 ;
        RECT 116.785 43.745 119.375 44.835 ;
        RECT 118.165 43.225 119.375 43.745 ;
        RECT 120.005 43.670 120.295 44.835 ;
        RECT 120.465 44.400 125.810 44.835 ;
        RECT 125.985 44.400 131.330 44.835 ;
        RECT 131.505 44.400 136.850 44.835 ;
        RECT 137.025 44.400 142.370 44.835 ;
        RECT 123.870 43.150 124.220 44.400 ;
        RECT 129.390 43.150 129.740 44.400 ;
        RECT 134.910 43.150 135.260 44.400 ;
        RECT 140.430 43.150 140.780 44.400 ;
        RECT 143.005 43.745 144.215 44.835 ;
        RECT 143.005 43.205 143.525 43.745 ;
        RECT 56.295 40.655 56.815 41.195 ;
        RECT 55.605 39.565 56.815 40.655 ;
        RECT 60.390 40.000 60.740 41.250 ;
        RECT 65.910 40.000 66.260 41.250 ;
        RECT 71.430 40.000 71.780 41.250 ;
        RECT 76.950 40.000 77.300 41.250 ;
        RECT 79.985 40.655 80.735 41.175 ;
        RECT 56.985 39.565 62.330 40.000 ;
        RECT 62.505 39.565 67.850 40.000 ;
        RECT 68.025 39.565 73.370 40.000 ;
        RECT 73.545 39.565 78.890 40.000 ;
        RECT 79.065 39.565 80.735 40.655 ;
        RECT 81.365 39.565 81.655 40.730 ;
        RECT 85.230 40.000 85.580 41.250 ;
        RECT 90.750 40.000 91.100 41.250 ;
        RECT 96.270 40.000 96.620 41.250 ;
        RECT 101.790 40.000 102.140 41.250 ;
        RECT 105.285 40.655 106.495 41.175 ;
        RECT 81.825 39.565 87.170 40.000 ;
        RECT 87.345 39.565 92.690 40.000 ;
        RECT 92.865 39.565 98.210 40.000 ;
        RECT 98.385 39.565 103.730 40.000 ;
        RECT 103.905 39.565 106.495 40.655 ;
        RECT 107.125 39.565 107.415 40.730 ;
        RECT 110.990 40.000 111.340 41.250 ;
        RECT 116.510 40.000 116.860 41.250 ;
        RECT 122.030 40.000 122.380 41.250 ;
        RECT 127.550 40.000 127.900 41.250 ;
        RECT 131.045 40.655 132.255 41.175 ;
        RECT 107.585 39.565 112.930 40.000 ;
        RECT 113.105 39.565 118.450 40.000 ;
        RECT 118.625 39.565 123.970 40.000 ;
        RECT 124.145 39.565 129.490 40.000 ;
        RECT 129.665 39.565 132.255 40.655 ;
        RECT 132.885 39.565 133.175 40.730 ;
        RECT 136.750 40.000 137.100 41.250 ;
        RECT 140.685 40.655 142.375 41.175 ;
        RECT 133.345 39.565 138.690 40.000 ;
        RECT 138.865 39.565 142.375 40.655 ;
        RECT 143.005 40.655 143.525 41.195 ;
        RECT 143.005 39.565 144.215 40.655 ;
        RECT 55.520 39.395 144.300 39.565 ;
        RECT 55.605 38.305 56.815 39.395 ;
        RECT 56.985 38.960 62.330 39.395 ;
        RECT 62.505 38.960 67.850 39.395 ;
        RECT 56.295 37.765 56.815 38.305 ;
        RECT 60.390 37.710 60.740 38.960 ;
        RECT 65.910 37.710 66.260 38.960 ;
        RECT 68.485 38.230 68.775 39.395 ;
        RECT 68.945 38.960 74.290 39.395 ;
        RECT 74.465 38.960 79.810 39.395 ;
        RECT 79.985 38.960 85.330 39.395 ;
        RECT 85.505 38.960 90.850 39.395 ;
        RECT 72.350 37.710 72.700 38.960 ;
        RECT 77.870 37.710 78.220 38.960 ;
        RECT 83.390 37.710 83.740 38.960 ;
        RECT 88.910 37.710 89.260 38.960 ;
        RECT 91.025 38.305 93.615 39.395 ;
        RECT 92.405 37.785 93.615 38.305 ;
        RECT 94.245 38.230 94.535 39.395 ;
        RECT 94.705 38.960 100.050 39.395 ;
        RECT 100.225 38.960 105.570 39.395 ;
        RECT 105.745 38.960 111.090 39.395 ;
        RECT 111.265 38.960 116.610 39.395 ;
        RECT 98.110 37.710 98.460 38.960 ;
        RECT 103.630 37.710 103.980 38.960 ;
        RECT 109.150 37.710 109.500 38.960 ;
        RECT 114.670 37.710 115.020 38.960 ;
        RECT 116.785 38.305 119.375 39.395 ;
        RECT 118.165 37.785 119.375 38.305 ;
        RECT 120.005 38.230 120.295 39.395 ;
        RECT 120.465 38.960 125.810 39.395 ;
        RECT 125.985 38.960 131.330 39.395 ;
        RECT 131.505 38.960 136.850 39.395 ;
        RECT 137.025 38.960 142.370 39.395 ;
        RECT 123.870 37.710 124.220 38.960 ;
        RECT 129.390 37.710 129.740 38.960 ;
        RECT 134.910 37.710 135.260 38.960 ;
        RECT 140.430 37.710 140.780 38.960 ;
        RECT 143.005 38.305 144.215 39.395 ;
        RECT 143.005 37.765 143.525 38.305 ;
        RECT 56.295 35.215 56.815 35.755 ;
        RECT 55.605 34.125 56.815 35.215 ;
        RECT 60.390 34.560 60.740 35.810 ;
        RECT 65.910 34.560 66.260 35.810 ;
        RECT 71.430 34.560 71.780 35.810 ;
        RECT 76.950 34.560 77.300 35.810 ;
        RECT 79.985 35.215 80.735 35.735 ;
        RECT 56.985 34.125 62.330 34.560 ;
        RECT 62.505 34.125 67.850 34.560 ;
        RECT 68.025 34.125 73.370 34.560 ;
        RECT 73.545 34.125 78.890 34.560 ;
        RECT 79.065 34.125 80.735 35.215 ;
        RECT 81.365 34.125 81.655 35.290 ;
        RECT 85.230 34.560 85.580 35.810 ;
        RECT 90.750 34.560 91.100 35.810 ;
        RECT 96.270 34.560 96.620 35.810 ;
        RECT 101.790 34.560 102.140 35.810 ;
        RECT 105.285 35.215 106.495 35.735 ;
        RECT 81.825 34.125 87.170 34.560 ;
        RECT 87.345 34.125 92.690 34.560 ;
        RECT 92.865 34.125 98.210 34.560 ;
        RECT 98.385 34.125 103.730 34.560 ;
        RECT 103.905 34.125 106.495 35.215 ;
        RECT 107.125 34.125 107.415 35.290 ;
        RECT 110.990 34.560 111.340 35.810 ;
        RECT 116.510 34.560 116.860 35.810 ;
        RECT 122.030 34.560 122.380 35.810 ;
        RECT 127.550 34.560 127.900 35.810 ;
        RECT 131.045 35.215 132.255 35.735 ;
        RECT 107.585 34.125 112.930 34.560 ;
        RECT 113.105 34.125 118.450 34.560 ;
        RECT 118.625 34.125 123.970 34.560 ;
        RECT 124.145 34.125 129.490 34.560 ;
        RECT 129.665 34.125 132.255 35.215 ;
        RECT 132.885 34.125 133.175 35.290 ;
        RECT 136.750 34.560 137.100 35.810 ;
        RECT 140.685 35.215 142.375 35.735 ;
        RECT 133.345 34.125 138.690 34.560 ;
        RECT 138.865 34.125 142.375 35.215 ;
        RECT 143.005 35.215 143.525 35.755 ;
        RECT 143.005 34.125 144.215 35.215 ;
        RECT 55.520 33.955 144.300 34.125 ;
        RECT 55.605 32.865 56.815 33.955 ;
        RECT 56.985 33.520 62.330 33.955 ;
        RECT 62.505 33.520 67.850 33.955 ;
        RECT 56.295 32.325 56.815 32.865 ;
        RECT 60.390 32.270 60.740 33.520 ;
        RECT 65.910 32.270 66.260 33.520 ;
        RECT 68.485 32.790 68.775 33.955 ;
        RECT 68.945 33.520 74.290 33.955 ;
        RECT 74.465 33.520 79.810 33.955 ;
        RECT 79.985 33.520 85.330 33.955 ;
        RECT 85.505 33.520 90.850 33.955 ;
        RECT 72.350 32.270 72.700 33.520 ;
        RECT 77.870 32.270 78.220 33.520 ;
        RECT 83.390 32.270 83.740 33.520 ;
        RECT 88.910 32.270 89.260 33.520 ;
        RECT 91.025 32.865 93.615 33.955 ;
        RECT 92.405 32.345 93.615 32.865 ;
        RECT 94.245 32.790 94.535 33.955 ;
        RECT 94.705 33.520 100.050 33.955 ;
        RECT 100.225 33.520 105.570 33.955 ;
        RECT 105.745 33.520 111.090 33.955 ;
        RECT 111.265 33.520 116.610 33.955 ;
        RECT 98.110 32.270 98.460 33.520 ;
        RECT 103.630 32.270 103.980 33.520 ;
        RECT 109.150 32.270 109.500 33.520 ;
        RECT 114.670 32.270 115.020 33.520 ;
        RECT 116.785 32.865 119.375 33.955 ;
        RECT 118.165 32.345 119.375 32.865 ;
        RECT 120.005 32.790 120.295 33.955 ;
        RECT 120.465 33.520 125.810 33.955 ;
        RECT 125.985 33.520 131.330 33.955 ;
        RECT 131.505 33.520 136.850 33.955 ;
        RECT 137.025 33.520 142.370 33.955 ;
        RECT 123.870 32.270 124.220 33.520 ;
        RECT 129.390 32.270 129.740 33.520 ;
        RECT 134.910 32.270 135.260 33.520 ;
        RECT 140.430 32.270 140.780 33.520 ;
        RECT 143.005 32.865 144.215 33.955 ;
        RECT 143.005 32.325 143.525 32.865 ;
        RECT 56.295 29.775 56.815 30.315 ;
        RECT 55.605 28.685 56.815 29.775 ;
        RECT 60.390 29.120 60.740 30.370 ;
        RECT 65.910 29.120 66.260 30.370 ;
        RECT 71.430 29.120 71.780 30.370 ;
        RECT 76.950 29.120 77.300 30.370 ;
        RECT 79.985 29.775 80.735 30.295 ;
        RECT 56.985 28.685 62.330 29.120 ;
        RECT 62.505 28.685 67.850 29.120 ;
        RECT 68.025 28.685 73.370 29.120 ;
        RECT 73.545 28.685 78.890 29.120 ;
        RECT 79.065 28.685 80.735 29.775 ;
        RECT 81.365 28.685 81.655 29.850 ;
        RECT 85.230 29.120 85.580 30.370 ;
        RECT 90.750 29.120 91.100 30.370 ;
        RECT 96.270 29.120 96.620 30.370 ;
        RECT 101.790 29.120 102.140 30.370 ;
        RECT 105.285 29.775 106.495 30.295 ;
        RECT 81.825 28.685 87.170 29.120 ;
        RECT 87.345 28.685 92.690 29.120 ;
        RECT 92.865 28.685 98.210 29.120 ;
        RECT 98.385 28.685 103.730 29.120 ;
        RECT 103.905 28.685 106.495 29.775 ;
        RECT 107.125 28.685 107.415 29.850 ;
        RECT 110.990 29.120 111.340 30.370 ;
        RECT 116.510 29.120 116.860 30.370 ;
        RECT 122.030 29.120 122.380 30.370 ;
        RECT 127.550 29.120 127.900 30.370 ;
        RECT 131.045 29.775 132.255 30.295 ;
        RECT 107.585 28.685 112.930 29.120 ;
        RECT 113.105 28.685 118.450 29.120 ;
        RECT 118.625 28.685 123.970 29.120 ;
        RECT 124.145 28.685 129.490 29.120 ;
        RECT 129.665 28.685 132.255 29.775 ;
        RECT 132.885 28.685 133.175 29.850 ;
        RECT 136.750 29.120 137.100 30.370 ;
        RECT 140.685 29.775 142.375 30.295 ;
        RECT 133.345 28.685 138.690 29.120 ;
        RECT 138.865 28.685 142.375 29.775 ;
        RECT 143.005 29.775 143.525 30.315 ;
        RECT 143.005 28.685 144.215 29.775 ;
        RECT 55.520 28.515 144.300 28.685 ;
        RECT 55.605 27.425 56.815 28.515 ;
        RECT 56.985 28.080 62.330 28.515 ;
        RECT 62.505 28.080 67.850 28.515 ;
        RECT 56.295 26.885 56.815 27.425 ;
        RECT 60.390 26.830 60.740 28.080 ;
        RECT 65.910 26.830 66.260 28.080 ;
        RECT 68.485 27.350 68.775 28.515 ;
        RECT 68.945 28.080 74.290 28.515 ;
        RECT 74.465 28.080 79.810 28.515 ;
        RECT 72.350 26.830 72.700 28.080 ;
        RECT 77.870 26.830 78.220 28.080 ;
        RECT 79.985 27.425 81.195 28.515 ;
        RECT 80.675 26.885 81.195 27.425 ;
        RECT 81.365 27.350 81.655 28.515 ;
        RECT 81.825 28.080 87.170 28.515 ;
        RECT 87.345 28.080 92.690 28.515 ;
        RECT 85.230 26.830 85.580 28.080 ;
        RECT 90.750 26.830 91.100 28.080 ;
        RECT 92.865 27.425 94.075 28.515 ;
        RECT 93.555 26.885 94.075 27.425 ;
        RECT 94.245 27.350 94.535 28.515 ;
        RECT 94.705 28.080 100.050 28.515 ;
        RECT 100.225 28.080 105.570 28.515 ;
        RECT 98.110 26.830 98.460 28.080 ;
        RECT 103.630 26.830 103.980 28.080 ;
        RECT 105.745 27.425 106.955 28.515 ;
        RECT 106.435 26.885 106.955 27.425 ;
        RECT 107.125 27.350 107.415 28.515 ;
        RECT 107.585 28.080 112.930 28.515 ;
        RECT 113.105 28.080 118.450 28.515 ;
        RECT 110.990 26.830 111.340 28.080 ;
        RECT 116.510 26.830 116.860 28.080 ;
        RECT 118.625 27.425 119.835 28.515 ;
        RECT 119.315 26.885 119.835 27.425 ;
        RECT 120.005 27.350 120.295 28.515 ;
        RECT 120.465 28.080 125.810 28.515 ;
        RECT 125.985 28.080 131.330 28.515 ;
        RECT 123.870 26.830 124.220 28.080 ;
        RECT 129.390 26.830 129.740 28.080 ;
        RECT 131.505 27.425 132.715 28.515 ;
        RECT 132.195 26.885 132.715 27.425 ;
        RECT 132.885 27.350 133.175 28.515 ;
        RECT 133.345 28.080 138.690 28.515 ;
        RECT 136.750 26.830 137.100 28.080 ;
        RECT 138.865 27.425 142.375 28.515 ;
        RECT 140.685 26.905 142.375 27.425 ;
        RECT 143.005 27.425 144.215 28.515 ;
        RECT 143.005 26.885 143.525 27.425 ;
      LAYER mcon ;
        RECT 55.665 99.235 55.835 99.405 ;
        RECT 56.125 99.235 56.295 99.405 ;
        RECT 56.585 99.235 56.755 99.405 ;
        RECT 57.045 99.235 57.215 99.405 ;
        RECT 57.505 99.235 57.675 99.405 ;
        RECT 57.965 99.235 58.135 99.405 ;
        RECT 58.425 99.235 58.595 99.405 ;
        RECT 58.885 99.235 59.055 99.405 ;
        RECT 59.345 99.235 59.515 99.405 ;
        RECT 59.805 99.235 59.975 99.405 ;
        RECT 60.265 99.235 60.435 99.405 ;
        RECT 60.725 99.235 60.895 99.405 ;
        RECT 61.185 99.235 61.355 99.405 ;
        RECT 61.645 99.235 61.815 99.405 ;
        RECT 62.105 99.235 62.275 99.405 ;
        RECT 62.565 99.235 62.735 99.405 ;
        RECT 63.025 99.235 63.195 99.405 ;
        RECT 63.485 99.235 63.655 99.405 ;
        RECT 63.945 99.235 64.115 99.405 ;
        RECT 64.405 99.235 64.575 99.405 ;
        RECT 64.865 99.235 65.035 99.405 ;
        RECT 65.325 99.235 65.495 99.405 ;
        RECT 65.785 99.235 65.955 99.405 ;
        RECT 66.245 99.235 66.415 99.405 ;
        RECT 66.705 99.235 66.875 99.405 ;
        RECT 67.165 99.235 67.335 99.405 ;
        RECT 67.625 99.235 67.795 99.405 ;
        RECT 68.085 99.235 68.255 99.405 ;
        RECT 68.545 99.235 68.715 99.405 ;
        RECT 69.005 99.235 69.175 99.405 ;
        RECT 69.465 99.235 69.635 99.405 ;
        RECT 69.925 99.235 70.095 99.405 ;
        RECT 70.385 99.235 70.555 99.405 ;
        RECT 70.845 99.235 71.015 99.405 ;
        RECT 71.305 99.235 71.475 99.405 ;
        RECT 71.765 99.235 71.935 99.405 ;
        RECT 72.225 99.235 72.395 99.405 ;
        RECT 72.685 99.235 72.855 99.405 ;
        RECT 73.145 99.235 73.315 99.405 ;
        RECT 73.605 99.235 73.775 99.405 ;
        RECT 74.065 99.235 74.235 99.405 ;
        RECT 74.525 99.235 74.695 99.405 ;
        RECT 74.985 99.235 75.155 99.405 ;
        RECT 75.445 99.235 75.615 99.405 ;
        RECT 75.905 99.235 76.075 99.405 ;
        RECT 76.365 99.235 76.535 99.405 ;
        RECT 76.825 99.235 76.995 99.405 ;
        RECT 77.285 99.235 77.455 99.405 ;
        RECT 77.745 99.235 77.915 99.405 ;
        RECT 78.205 99.235 78.375 99.405 ;
        RECT 78.665 99.235 78.835 99.405 ;
        RECT 79.125 99.235 79.295 99.405 ;
        RECT 79.585 99.235 79.755 99.405 ;
        RECT 80.045 99.235 80.215 99.405 ;
        RECT 80.505 99.235 80.675 99.405 ;
        RECT 80.965 99.235 81.135 99.405 ;
        RECT 81.425 99.235 81.595 99.405 ;
        RECT 81.885 99.235 82.055 99.405 ;
        RECT 82.345 99.235 82.515 99.405 ;
        RECT 82.805 99.235 82.975 99.405 ;
        RECT 83.265 99.235 83.435 99.405 ;
        RECT 83.725 99.235 83.895 99.405 ;
        RECT 84.185 99.235 84.355 99.405 ;
        RECT 84.645 99.235 84.815 99.405 ;
        RECT 85.105 99.235 85.275 99.405 ;
        RECT 85.565 99.235 85.735 99.405 ;
        RECT 86.025 99.235 86.195 99.405 ;
        RECT 86.485 99.235 86.655 99.405 ;
        RECT 86.945 99.235 87.115 99.405 ;
        RECT 87.405 99.235 87.575 99.405 ;
        RECT 87.865 99.235 88.035 99.405 ;
        RECT 88.325 99.235 88.495 99.405 ;
        RECT 88.785 99.235 88.955 99.405 ;
        RECT 89.245 99.235 89.415 99.405 ;
        RECT 89.705 99.235 89.875 99.405 ;
        RECT 90.165 99.235 90.335 99.405 ;
        RECT 90.625 99.235 90.795 99.405 ;
        RECT 91.085 99.235 91.255 99.405 ;
        RECT 91.545 99.235 91.715 99.405 ;
        RECT 92.005 99.235 92.175 99.405 ;
        RECT 92.465 99.235 92.635 99.405 ;
        RECT 92.925 99.235 93.095 99.405 ;
        RECT 93.385 99.235 93.555 99.405 ;
        RECT 93.845 99.235 94.015 99.405 ;
        RECT 94.305 99.235 94.475 99.405 ;
        RECT 94.765 99.235 94.935 99.405 ;
        RECT 95.225 99.235 95.395 99.405 ;
        RECT 95.685 99.235 95.855 99.405 ;
        RECT 96.145 99.235 96.315 99.405 ;
        RECT 96.605 99.235 96.775 99.405 ;
        RECT 97.065 99.235 97.235 99.405 ;
        RECT 97.525 99.235 97.695 99.405 ;
        RECT 97.985 99.235 98.155 99.405 ;
        RECT 98.445 99.235 98.615 99.405 ;
        RECT 98.905 99.235 99.075 99.405 ;
        RECT 99.365 99.235 99.535 99.405 ;
        RECT 99.825 99.235 99.995 99.405 ;
        RECT 100.285 99.235 100.455 99.405 ;
        RECT 100.745 99.235 100.915 99.405 ;
        RECT 101.205 99.235 101.375 99.405 ;
        RECT 101.665 99.235 101.835 99.405 ;
        RECT 102.125 99.235 102.295 99.405 ;
        RECT 102.585 99.235 102.755 99.405 ;
        RECT 103.045 99.235 103.215 99.405 ;
        RECT 103.505 99.235 103.675 99.405 ;
        RECT 103.965 99.235 104.135 99.405 ;
        RECT 104.425 99.235 104.595 99.405 ;
        RECT 104.885 99.235 105.055 99.405 ;
        RECT 105.345 99.235 105.515 99.405 ;
        RECT 105.805 99.235 105.975 99.405 ;
        RECT 106.265 99.235 106.435 99.405 ;
        RECT 106.725 99.235 106.895 99.405 ;
        RECT 107.185 99.235 107.355 99.405 ;
        RECT 107.645 99.235 107.815 99.405 ;
        RECT 108.105 99.235 108.275 99.405 ;
        RECT 108.565 99.235 108.735 99.405 ;
        RECT 109.025 99.235 109.195 99.405 ;
        RECT 109.485 99.235 109.655 99.405 ;
        RECT 109.945 99.235 110.115 99.405 ;
        RECT 110.405 99.235 110.575 99.405 ;
        RECT 110.865 99.235 111.035 99.405 ;
        RECT 111.325 99.235 111.495 99.405 ;
        RECT 111.785 99.235 111.955 99.405 ;
        RECT 112.245 99.235 112.415 99.405 ;
        RECT 112.705 99.235 112.875 99.405 ;
        RECT 113.165 99.235 113.335 99.405 ;
        RECT 113.625 99.235 113.795 99.405 ;
        RECT 114.085 99.235 114.255 99.405 ;
        RECT 114.545 99.235 114.715 99.405 ;
        RECT 115.005 99.235 115.175 99.405 ;
        RECT 115.465 99.235 115.635 99.405 ;
        RECT 115.925 99.235 116.095 99.405 ;
        RECT 116.385 99.235 116.555 99.405 ;
        RECT 116.845 99.235 117.015 99.405 ;
        RECT 117.305 99.235 117.475 99.405 ;
        RECT 117.765 99.235 117.935 99.405 ;
        RECT 118.225 99.235 118.395 99.405 ;
        RECT 118.685 99.235 118.855 99.405 ;
        RECT 119.145 99.235 119.315 99.405 ;
        RECT 119.605 99.235 119.775 99.405 ;
        RECT 120.065 99.235 120.235 99.405 ;
        RECT 120.525 99.235 120.695 99.405 ;
        RECT 120.985 99.235 121.155 99.405 ;
        RECT 121.445 99.235 121.615 99.405 ;
        RECT 121.905 99.235 122.075 99.405 ;
        RECT 122.365 99.235 122.535 99.405 ;
        RECT 122.825 99.235 122.995 99.405 ;
        RECT 123.285 99.235 123.455 99.405 ;
        RECT 123.745 99.235 123.915 99.405 ;
        RECT 124.205 99.235 124.375 99.405 ;
        RECT 124.665 99.235 124.835 99.405 ;
        RECT 125.125 99.235 125.295 99.405 ;
        RECT 125.585 99.235 125.755 99.405 ;
        RECT 126.045 99.235 126.215 99.405 ;
        RECT 126.505 99.235 126.675 99.405 ;
        RECT 126.965 99.235 127.135 99.405 ;
        RECT 127.425 99.235 127.595 99.405 ;
        RECT 127.885 99.235 128.055 99.405 ;
        RECT 128.345 99.235 128.515 99.405 ;
        RECT 128.805 99.235 128.975 99.405 ;
        RECT 129.265 99.235 129.435 99.405 ;
        RECT 129.725 99.235 129.895 99.405 ;
        RECT 130.185 99.235 130.355 99.405 ;
        RECT 130.645 99.235 130.815 99.405 ;
        RECT 131.105 99.235 131.275 99.405 ;
        RECT 131.565 99.235 131.735 99.405 ;
        RECT 132.025 99.235 132.195 99.405 ;
        RECT 132.485 99.235 132.655 99.405 ;
        RECT 132.945 99.235 133.115 99.405 ;
        RECT 133.405 99.235 133.575 99.405 ;
        RECT 133.865 99.235 134.035 99.405 ;
        RECT 134.325 99.235 134.495 99.405 ;
        RECT 134.785 99.235 134.955 99.405 ;
        RECT 135.245 99.235 135.415 99.405 ;
        RECT 135.705 99.235 135.875 99.405 ;
        RECT 136.165 99.235 136.335 99.405 ;
        RECT 136.625 99.235 136.795 99.405 ;
        RECT 137.085 99.235 137.255 99.405 ;
        RECT 137.545 99.235 137.715 99.405 ;
        RECT 138.005 99.235 138.175 99.405 ;
        RECT 138.465 99.235 138.635 99.405 ;
        RECT 138.925 99.235 139.095 99.405 ;
        RECT 139.385 99.235 139.555 99.405 ;
        RECT 139.845 99.235 140.015 99.405 ;
        RECT 140.305 99.235 140.475 99.405 ;
        RECT 140.765 99.235 140.935 99.405 ;
        RECT 141.225 99.235 141.395 99.405 ;
        RECT 141.685 99.235 141.855 99.405 ;
        RECT 142.145 99.235 142.315 99.405 ;
        RECT 142.605 99.235 142.775 99.405 ;
        RECT 143.065 99.235 143.235 99.405 ;
        RECT 143.525 99.235 143.695 99.405 ;
        RECT 143.985 99.235 144.155 99.405 ;
        RECT 55.665 93.795 55.835 93.965 ;
        RECT 56.125 93.795 56.295 93.965 ;
        RECT 56.585 93.795 56.755 93.965 ;
        RECT 57.045 93.795 57.215 93.965 ;
        RECT 57.505 93.795 57.675 93.965 ;
        RECT 57.965 93.795 58.135 93.965 ;
        RECT 58.425 93.795 58.595 93.965 ;
        RECT 58.885 93.795 59.055 93.965 ;
        RECT 59.345 93.795 59.515 93.965 ;
        RECT 59.805 93.795 59.975 93.965 ;
        RECT 60.265 93.795 60.435 93.965 ;
        RECT 60.725 93.795 60.895 93.965 ;
        RECT 61.185 93.795 61.355 93.965 ;
        RECT 61.645 93.795 61.815 93.965 ;
        RECT 62.105 93.795 62.275 93.965 ;
        RECT 62.565 93.795 62.735 93.965 ;
        RECT 63.025 93.795 63.195 93.965 ;
        RECT 63.485 93.795 63.655 93.965 ;
        RECT 63.945 93.795 64.115 93.965 ;
        RECT 64.405 93.795 64.575 93.965 ;
        RECT 64.865 93.795 65.035 93.965 ;
        RECT 65.325 93.795 65.495 93.965 ;
        RECT 65.785 93.795 65.955 93.965 ;
        RECT 66.245 93.795 66.415 93.965 ;
        RECT 66.705 93.795 66.875 93.965 ;
        RECT 67.165 93.795 67.335 93.965 ;
        RECT 67.625 93.795 67.795 93.965 ;
        RECT 68.085 93.795 68.255 93.965 ;
        RECT 68.545 93.795 68.715 93.965 ;
        RECT 69.005 93.795 69.175 93.965 ;
        RECT 69.465 93.795 69.635 93.965 ;
        RECT 69.925 93.795 70.095 93.965 ;
        RECT 70.385 93.795 70.555 93.965 ;
        RECT 70.845 93.795 71.015 93.965 ;
        RECT 71.305 93.795 71.475 93.965 ;
        RECT 71.765 93.795 71.935 93.965 ;
        RECT 72.225 93.795 72.395 93.965 ;
        RECT 72.685 93.795 72.855 93.965 ;
        RECT 73.145 93.795 73.315 93.965 ;
        RECT 73.605 93.795 73.775 93.965 ;
        RECT 74.065 93.795 74.235 93.965 ;
        RECT 74.525 93.795 74.695 93.965 ;
        RECT 74.985 93.795 75.155 93.965 ;
        RECT 75.445 93.795 75.615 93.965 ;
        RECT 75.905 93.795 76.075 93.965 ;
        RECT 76.365 93.795 76.535 93.965 ;
        RECT 76.825 93.795 76.995 93.965 ;
        RECT 77.285 93.795 77.455 93.965 ;
        RECT 77.745 93.795 77.915 93.965 ;
        RECT 78.205 93.795 78.375 93.965 ;
        RECT 78.665 93.795 78.835 93.965 ;
        RECT 79.125 93.795 79.295 93.965 ;
        RECT 79.585 93.795 79.755 93.965 ;
        RECT 80.045 93.795 80.215 93.965 ;
        RECT 80.505 93.795 80.675 93.965 ;
        RECT 80.965 93.795 81.135 93.965 ;
        RECT 81.425 93.795 81.595 93.965 ;
        RECT 81.885 93.795 82.055 93.965 ;
        RECT 82.345 93.795 82.515 93.965 ;
        RECT 82.805 93.795 82.975 93.965 ;
        RECT 83.265 93.795 83.435 93.965 ;
        RECT 83.725 93.795 83.895 93.965 ;
        RECT 84.185 93.795 84.355 93.965 ;
        RECT 84.645 93.795 84.815 93.965 ;
        RECT 85.105 93.795 85.275 93.965 ;
        RECT 85.565 93.795 85.735 93.965 ;
        RECT 86.025 93.795 86.195 93.965 ;
        RECT 86.485 93.795 86.655 93.965 ;
        RECT 86.945 93.795 87.115 93.965 ;
        RECT 87.405 93.795 87.575 93.965 ;
        RECT 87.865 93.795 88.035 93.965 ;
        RECT 88.325 93.795 88.495 93.965 ;
        RECT 88.785 93.795 88.955 93.965 ;
        RECT 89.245 93.795 89.415 93.965 ;
        RECT 89.705 93.795 89.875 93.965 ;
        RECT 90.165 93.795 90.335 93.965 ;
        RECT 90.625 93.795 90.795 93.965 ;
        RECT 91.085 93.795 91.255 93.965 ;
        RECT 91.545 93.795 91.715 93.965 ;
        RECT 92.005 93.795 92.175 93.965 ;
        RECT 92.465 93.795 92.635 93.965 ;
        RECT 92.925 93.795 93.095 93.965 ;
        RECT 93.385 93.795 93.555 93.965 ;
        RECT 93.845 93.795 94.015 93.965 ;
        RECT 94.305 93.795 94.475 93.965 ;
        RECT 94.765 93.795 94.935 93.965 ;
        RECT 95.225 93.795 95.395 93.965 ;
        RECT 95.685 93.795 95.855 93.965 ;
        RECT 96.145 93.795 96.315 93.965 ;
        RECT 96.605 93.795 96.775 93.965 ;
        RECT 97.065 93.795 97.235 93.965 ;
        RECT 97.525 93.795 97.695 93.965 ;
        RECT 97.985 93.795 98.155 93.965 ;
        RECT 98.445 93.795 98.615 93.965 ;
        RECT 98.905 93.795 99.075 93.965 ;
        RECT 99.365 93.795 99.535 93.965 ;
        RECT 99.825 93.795 99.995 93.965 ;
        RECT 100.285 93.795 100.455 93.965 ;
        RECT 100.745 93.795 100.915 93.965 ;
        RECT 101.205 93.795 101.375 93.965 ;
        RECT 101.665 93.795 101.835 93.965 ;
        RECT 102.125 93.795 102.295 93.965 ;
        RECT 102.585 93.795 102.755 93.965 ;
        RECT 103.045 93.795 103.215 93.965 ;
        RECT 103.505 93.795 103.675 93.965 ;
        RECT 103.965 93.795 104.135 93.965 ;
        RECT 104.425 93.795 104.595 93.965 ;
        RECT 104.885 93.795 105.055 93.965 ;
        RECT 105.345 93.795 105.515 93.965 ;
        RECT 105.805 93.795 105.975 93.965 ;
        RECT 106.265 93.795 106.435 93.965 ;
        RECT 106.725 93.795 106.895 93.965 ;
        RECT 107.185 93.795 107.355 93.965 ;
        RECT 107.645 93.795 107.815 93.965 ;
        RECT 108.105 93.795 108.275 93.965 ;
        RECT 108.565 93.795 108.735 93.965 ;
        RECT 109.025 93.795 109.195 93.965 ;
        RECT 109.485 93.795 109.655 93.965 ;
        RECT 109.945 93.795 110.115 93.965 ;
        RECT 110.405 93.795 110.575 93.965 ;
        RECT 110.865 93.795 111.035 93.965 ;
        RECT 111.325 93.795 111.495 93.965 ;
        RECT 111.785 93.795 111.955 93.965 ;
        RECT 112.245 93.795 112.415 93.965 ;
        RECT 112.705 93.795 112.875 93.965 ;
        RECT 113.165 93.795 113.335 93.965 ;
        RECT 113.625 93.795 113.795 93.965 ;
        RECT 114.085 93.795 114.255 93.965 ;
        RECT 114.545 93.795 114.715 93.965 ;
        RECT 115.005 93.795 115.175 93.965 ;
        RECT 115.465 93.795 115.635 93.965 ;
        RECT 115.925 93.795 116.095 93.965 ;
        RECT 116.385 93.795 116.555 93.965 ;
        RECT 116.845 93.795 117.015 93.965 ;
        RECT 117.305 93.795 117.475 93.965 ;
        RECT 117.765 93.795 117.935 93.965 ;
        RECT 118.225 93.795 118.395 93.965 ;
        RECT 118.685 93.795 118.855 93.965 ;
        RECT 119.145 93.795 119.315 93.965 ;
        RECT 119.605 93.795 119.775 93.965 ;
        RECT 120.065 93.795 120.235 93.965 ;
        RECT 120.525 93.795 120.695 93.965 ;
        RECT 120.985 93.795 121.155 93.965 ;
        RECT 121.445 93.795 121.615 93.965 ;
        RECT 121.905 93.795 122.075 93.965 ;
        RECT 122.365 93.795 122.535 93.965 ;
        RECT 122.825 93.795 122.995 93.965 ;
        RECT 123.285 93.795 123.455 93.965 ;
        RECT 123.745 93.795 123.915 93.965 ;
        RECT 124.205 93.795 124.375 93.965 ;
        RECT 124.665 93.795 124.835 93.965 ;
        RECT 125.125 93.795 125.295 93.965 ;
        RECT 125.585 93.795 125.755 93.965 ;
        RECT 126.045 93.795 126.215 93.965 ;
        RECT 126.505 93.795 126.675 93.965 ;
        RECT 126.965 93.795 127.135 93.965 ;
        RECT 127.425 93.795 127.595 93.965 ;
        RECT 127.885 93.795 128.055 93.965 ;
        RECT 128.345 93.795 128.515 93.965 ;
        RECT 128.805 93.795 128.975 93.965 ;
        RECT 129.265 93.795 129.435 93.965 ;
        RECT 129.725 93.795 129.895 93.965 ;
        RECT 130.185 93.795 130.355 93.965 ;
        RECT 130.645 93.795 130.815 93.965 ;
        RECT 131.105 93.795 131.275 93.965 ;
        RECT 131.565 93.795 131.735 93.965 ;
        RECT 132.025 93.795 132.195 93.965 ;
        RECT 132.485 93.795 132.655 93.965 ;
        RECT 132.945 93.795 133.115 93.965 ;
        RECT 133.405 93.795 133.575 93.965 ;
        RECT 133.865 93.795 134.035 93.965 ;
        RECT 134.325 93.795 134.495 93.965 ;
        RECT 134.785 93.795 134.955 93.965 ;
        RECT 135.245 93.795 135.415 93.965 ;
        RECT 135.705 93.795 135.875 93.965 ;
        RECT 136.165 93.795 136.335 93.965 ;
        RECT 136.625 93.795 136.795 93.965 ;
        RECT 137.085 93.795 137.255 93.965 ;
        RECT 137.545 93.795 137.715 93.965 ;
        RECT 138.005 93.795 138.175 93.965 ;
        RECT 138.465 93.795 138.635 93.965 ;
        RECT 138.925 93.795 139.095 93.965 ;
        RECT 139.385 93.795 139.555 93.965 ;
        RECT 139.845 93.795 140.015 93.965 ;
        RECT 140.305 93.795 140.475 93.965 ;
        RECT 140.765 93.795 140.935 93.965 ;
        RECT 141.225 93.795 141.395 93.965 ;
        RECT 141.685 93.795 141.855 93.965 ;
        RECT 142.145 93.795 142.315 93.965 ;
        RECT 142.605 93.795 142.775 93.965 ;
        RECT 143.065 93.795 143.235 93.965 ;
        RECT 143.525 93.795 143.695 93.965 ;
        RECT 143.985 93.795 144.155 93.965 ;
        RECT 55.665 88.355 55.835 88.525 ;
        RECT 56.125 88.355 56.295 88.525 ;
        RECT 56.585 88.355 56.755 88.525 ;
        RECT 57.045 88.355 57.215 88.525 ;
        RECT 57.505 88.355 57.675 88.525 ;
        RECT 57.965 88.355 58.135 88.525 ;
        RECT 58.425 88.355 58.595 88.525 ;
        RECT 58.885 88.355 59.055 88.525 ;
        RECT 59.345 88.355 59.515 88.525 ;
        RECT 59.805 88.355 59.975 88.525 ;
        RECT 60.265 88.355 60.435 88.525 ;
        RECT 60.725 88.355 60.895 88.525 ;
        RECT 61.185 88.355 61.355 88.525 ;
        RECT 61.645 88.355 61.815 88.525 ;
        RECT 62.105 88.355 62.275 88.525 ;
        RECT 62.565 88.355 62.735 88.525 ;
        RECT 63.025 88.355 63.195 88.525 ;
        RECT 63.485 88.355 63.655 88.525 ;
        RECT 63.945 88.355 64.115 88.525 ;
        RECT 64.405 88.355 64.575 88.525 ;
        RECT 64.865 88.355 65.035 88.525 ;
        RECT 65.325 88.355 65.495 88.525 ;
        RECT 65.785 88.355 65.955 88.525 ;
        RECT 66.245 88.355 66.415 88.525 ;
        RECT 66.705 88.355 66.875 88.525 ;
        RECT 67.165 88.355 67.335 88.525 ;
        RECT 67.625 88.355 67.795 88.525 ;
        RECT 68.085 88.355 68.255 88.525 ;
        RECT 68.545 88.355 68.715 88.525 ;
        RECT 69.005 88.355 69.175 88.525 ;
        RECT 69.465 88.355 69.635 88.525 ;
        RECT 69.925 88.355 70.095 88.525 ;
        RECT 70.385 88.355 70.555 88.525 ;
        RECT 70.845 88.355 71.015 88.525 ;
        RECT 71.305 88.355 71.475 88.525 ;
        RECT 71.765 88.355 71.935 88.525 ;
        RECT 72.225 88.355 72.395 88.525 ;
        RECT 72.685 88.355 72.855 88.525 ;
        RECT 73.145 88.355 73.315 88.525 ;
        RECT 73.605 88.355 73.775 88.525 ;
        RECT 74.065 88.355 74.235 88.525 ;
        RECT 74.525 88.355 74.695 88.525 ;
        RECT 74.985 88.355 75.155 88.525 ;
        RECT 75.445 88.355 75.615 88.525 ;
        RECT 75.905 88.355 76.075 88.525 ;
        RECT 76.365 88.355 76.535 88.525 ;
        RECT 76.825 88.355 76.995 88.525 ;
        RECT 77.285 88.355 77.455 88.525 ;
        RECT 77.745 88.355 77.915 88.525 ;
        RECT 78.205 88.355 78.375 88.525 ;
        RECT 78.665 88.355 78.835 88.525 ;
        RECT 79.125 88.355 79.295 88.525 ;
        RECT 79.585 88.355 79.755 88.525 ;
        RECT 80.045 88.355 80.215 88.525 ;
        RECT 80.505 88.355 80.675 88.525 ;
        RECT 80.965 88.355 81.135 88.525 ;
        RECT 81.425 88.355 81.595 88.525 ;
        RECT 81.885 88.355 82.055 88.525 ;
        RECT 82.345 88.355 82.515 88.525 ;
        RECT 82.805 88.355 82.975 88.525 ;
        RECT 83.265 88.355 83.435 88.525 ;
        RECT 83.725 88.355 83.895 88.525 ;
        RECT 84.185 88.355 84.355 88.525 ;
        RECT 84.645 88.355 84.815 88.525 ;
        RECT 85.105 88.355 85.275 88.525 ;
        RECT 85.565 88.355 85.735 88.525 ;
        RECT 86.025 88.355 86.195 88.525 ;
        RECT 86.485 88.355 86.655 88.525 ;
        RECT 86.945 88.355 87.115 88.525 ;
        RECT 87.405 88.355 87.575 88.525 ;
        RECT 87.865 88.355 88.035 88.525 ;
        RECT 88.325 88.355 88.495 88.525 ;
        RECT 88.785 88.355 88.955 88.525 ;
        RECT 89.245 88.355 89.415 88.525 ;
        RECT 89.705 88.355 89.875 88.525 ;
        RECT 90.165 88.355 90.335 88.525 ;
        RECT 90.625 88.355 90.795 88.525 ;
        RECT 91.085 88.355 91.255 88.525 ;
        RECT 91.545 88.355 91.715 88.525 ;
        RECT 92.005 88.355 92.175 88.525 ;
        RECT 92.465 88.355 92.635 88.525 ;
        RECT 92.925 88.355 93.095 88.525 ;
        RECT 93.385 88.355 93.555 88.525 ;
        RECT 93.845 88.355 94.015 88.525 ;
        RECT 94.305 88.355 94.475 88.525 ;
        RECT 94.765 88.355 94.935 88.525 ;
        RECT 95.225 88.355 95.395 88.525 ;
        RECT 95.685 88.355 95.855 88.525 ;
        RECT 96.145 88.355 96.315 88.525 ;
        RECT 96.605 88.355 96.775 88.525 ;
        RECT 97.065 88.355 97.235 88.525 ;
        RECT 97.525 88.355 97.695 88.525 ;
        RECT 97.985 88.355 98.155 88.525 ;
        RECT 98.445 88.355 98.615 88.525 ;
        RECT 98.905 88.355 99.075 88.525 ;
        RECT 99.365 88.355 99.535 88.525 ;
        RECT 99.825 88.355 99.995 88.525 ;
        RECT 100.285 88.355 100.455 88.525 ;
        RECT 100.745 88.355 100.915 88.525 ;
        RECT 101.205 88.355 101.375 88.525 ;
        RECT 101.665 88.355 101.835 88.525 ;
        RECT 102.125 88.355 102.295 88.525 ;
        RECT 102.585 88.355 102.755 88.525 ;
        RECT 103.045 88.355 103.215 88.525 ;
        RECT 103.505 88.355 103.675 88.525 ;
        RECT 103.965 88.355 104.135 88.525 ;
        RECT 104.425 88.355 104.595 88.525 ;
        RECT 104.885 88.355 105.055 88.525 ;
        RECT 105.345 88.355 105.515 88.525 ;
        RECT 105.805 88.355 105.975 88.525 ;
        RECT 106.265 88.355 106.435 88.525 ;
        RECT 106.725 88.355 106.895 88.525 ;
        RECT 107.185 88.355 107.355 88.525 ;
        RECT 107.645 88.355 107.815 88.525 ;
        RECT 108.105 88.355 108.275 88.525 ;
        RECT 108.565 88.355 108.735 88.525 ;
        RECT 109.025 88.355 109.195 88.525 ;
        RECT 109.485 88.355 109.655 88.525 ;
        RECT 109.945 88.355 110.115 88.525 ;
        RECT 110.405 88.355 110.575 88.525 ;
        RECT 110.865 88.355 111.035 88.525 ;
        RECT 111.325 88.355 111.495 88.525 ;
        RECT 111.785 88.355 111.955 88.525 ;
        RECT 112.245 88.355 112.415 88.525 ;
        RECT 112.705 88.355 112.875 88.525 ;
        RECT 113.165 88.355 113.335 88.525 ;
        RECT 113.625 88.355 113.795 88.525 ;
        RECT 114.085 88.355 114.255 88.525 ;
        RECT 114.545 88.355 114.715 88.525 ;
        RECT 115.005 88.355 115.175 88.525 ;
        RECT 115.465 88.355 115.635 88.525 ;
        RECT 115.925 88.355 116.095 88.525 ;
        RECT 116.385 88.355 116.555 88.525 ;
        RECT 116.845 88.355 117.015 88.525 ;
        RECT 117.305 88.355 117.475 88.525 ;
        RECT 117.765 88.355 117.935 88.525 ;
        RECT 118.225 88.355 118.395 88.525 ;
        RECT 118.685 88.355 118.855 88.525 ;
        RECT 119.145 88.355 119.315 88.525 ;
        RECT 119.605 88.355 119.775 88.525 ;
        RECT 120.065 88.355 120.235 88.525 ;
        RECT 120.525 88.355 120.695 88.525 ;
        RECT 120.985 88.355 121.155 88.525 ;
        RECT 121.445 88.355 121.615 88.525 ;
        RECT 121.905 88.355 122.075 88.525 ;
        RECT 122.365 88.355 122.535 88.525 ;
        RECT 122.825 88.355 122.995 88.525 ;
        RECT 123.285 88.355 123.455 88.525 ;
        RECT 123.745 88.355 123.915 88.525 ;
        RECT 124.205 88.355 124.375 88.525 ;
        RECT 124.665 88.355 124.835 88.525 ;
        RECT 125.125 88.355 125.295 88.525 ;
        RECT 125.585 88.355 125.755 88.525 ;
        RECT 126.045 88.355 126.215 88.525 ;
        RECT 126.505 88.355 126.675 88.525 ;
        RECT 126.965 88.355 127.135 88.525 ;
        RECT 127.425 88.355 127.595 88.525 ;
        RECT 127.885 88.355 128.055 88.525 ;
        RECT 128.345 88.355 128.515 88.525 ;
        RECT 128.805 88.355 128.975 88.525 ;
        RECT 129.265 88.355 129.435 88.525 ;
        RECT 129.725 88.355 129.895 88.525 ;
        RECT 130.185 88.355 130.355 88.525 ;
        RECT 130.645 88.355 130.815 88.525 ;
        RECT 131.105 88.355 131.275 88.525 ;
        RECT 131.565 88.355 131.735 88.525 ;
        RECT 132.025 88.355 132.195 88.525 ;
        RECT 132.485 88.355 132.655 88.525 ;
        RECT 132.945 88.355 133.115 88.525 ;
        RECT 133.405 88.355 133.575 88.525 ;
        RECT 133.865 88.355 134.035 88.525 ;
        RECT 134.325 88.355 134.495 88.525 ;
        RECT 134.785 88.355 134.955 88.525 ;
        RECT 135.245 88.355 135.415 88.525 ;
        RECT 135.705 88.355 135.875 88.525 ;
        RECT 136.165 88.355 136.335 88.525 ;
        RECT 136.625 88.355 136.795 88.525 ;
        RECT 137.085 88.355 137.255 88.525 ;
        RECT 137.545 88.355 137.715 88.525 ;
        RECT 138.005 88.355 138.175 88.525 ;
        RECT 138.465 88.355 138.635 88.525 ;
        RECT 138.925 88.355 139.095 88.525 ;
        RECT 139.385 88.355 139.555 88.525 ;
        RECT 139.845 88.355 140.015 88.525 ;
        RECT 140.305 88.355 140.475 88.525 ;
        RECT 140.765 88.355 140.935 88.525 ;
        RECT 141.225 88.355 141.395 88.525 ;
        RECT 141.685 88.355 141.855 88.525 ;
        RECT 142.145 88.355 142.315 88.525 ;
        RECT 142.605 88.355 142.775 88.525 ;
        RECT 143.065 88.355 143.235 88.525 ;
        RECT 143.525 88.355 143.695 88.525 ;
        RECT 143.985 88.355 144.155 88.525 ;
        RECT 55.665 82.915 55.835 83.085 ;
        RECT 56.125 82.915 56.295 83.085 ;
        RECT 56.585 82.915 56.755 83.085 ;
        RECT 57.045 82.915 57.215 83.085 ;
        RECT 57.505 82.915 57.675 83.085 ;
        RECT 57.965 82.915 58.135 83.085 ;
        RECT 58.425 82.915 58.595 83.085 ;
        RECT 58.885 82.915 59.055 83.085 ;
        RECT 59.345 82.915 59.515 83.085 ;
        RECT 59.805 82.915 59.975 83.085 ;
        RECT 60.265 82.915 60.435 83.085 ;
        RECT 60.725 82.915 60.895 83.085 ;
        RECT 61.185 82.915 61.355 83.085 ;
        RECT 61.645 82.915 61.815 83.085 ;
        RECT 62.105 82.915 62.275 83.085 ;
        RECT 62.565 82.915 62.735 83.085 ;
        RECT 63.025 82.915 63.195 83.085 ;
        RECT 63.485 82.915 63.655 83.085 ;
        RECT 63.945 82.915 64.115 83.085 ;
        RECT 64.405 82.915 64.575 83.085 ;
        RECT 64.865 82.915 65.035 83.085 ;
        RECT 65.325 82.915 65.495 83.085 ;
        RECT 65.785 82.915 65.955 83.085 ;
        RECT 66.245 82.915 66.415 83.085 ;
        RECT 66.705 82.915 66.875 83.085 ;
        RECT 67.165 82.915 67.335 83.085 ;
        RECT 67.625 82.915 67.795 83.085 ;
        RECT 68.085 82.915 68.255 83.085 ;
        RECT 68.545 82.915 68.715 83.085 ;
        RECT 69.005 82.915 69.175 83.085 ;
        RECT 69.465 82.915 69.635 83.085 ;
        RECT 69.925 82.915 70.095 83.085 ;
        RECT 70.385 82.915 70.555 83.085 ;
        RECT 70.845 82.915 71.015 83.085 ;
        RECT 71.305 82.915 71.475 83.085 ;
        RECT 71.765 82.915 71.935 83.085 ;
        RECT 72.225 82.915 72.395 83.085 ;
        RECT 72.685 82.915 72.855 83.085 ;
        RECT 73.145 82.915 73.315 83.085 ;
        RECT 73.605 82.915 73.775 83.085 ;
        RECT 74.065 82.915 74.235 83.085 ;
        RECT 74.525 82.915 74.695 83.085 ;
        RECT 74.985 82.915 75.155 83.085 ;
        RECT 75.445 82.915 75.615 83.085 ;
        RECT 75.905 82.915 76.075 83.085 ;
        RECT 76.365 82.915 76.535 83.085 ;
        RECT 76.825 82.915 76.995 83.085 ;
        RECT 77.285 82.915 77.455 83.085 ;
        RECT 77.745 82.915 77.915 83.085 ;
        RECT 78.205 82.915 78.375 83.085 ;
        RECT 78.665 82.915 78.835 83.085 ;
        RECT 79.125 82.915 79.295 83.085 ;
        RECT 79.585 82.915 79.755 83.085 ;
        RECT 80.045 82.915 80.215 83.085 ;
        RECT 80.505 82.915 80.675 83.085 ;
        RECT 80.965 82.915 81.135 83.085 ;
        RECT 81.425 82.915 81.595 83.085 ;
        RECT 81.885 82.915 82.055 83.085 ;
        RECT 82.345 82.915 82.515 83.085 ;
        RECT 82.805 82.915 82.975 83.085 ;
        RECT 83.265 82.915 83.435 83.085 ;
        RECT 83.725 82.915 83.895 83.085 ;
        RECT 84.185 82.915 84.355 83.085 ;
        RECT 84.645 82.915 84.815 83.085 ;
        RECT 85.105 82.915 85.275 83.085 ;
        RECT 85.565 82.915 85.735 83.085 ;
        RECT 86.025 82.915 86.195 83.085 ;
        RECT 86.485 82.915 86.655 83.085 ;
        RECT 86.945 82.915 87.115 83.085 ;
        RECT 87.405 82.915 87.575 83.085 ;
        RECT 87.865 82.915 88.035 83.085 ;
        RECT 88.325 82.915 88.495 83.085 ;
        RECT 88.785 82.915 88.955 83.085 ;
        RECT 89.245 82.915 89.415 83.085 ;
        RECT 89.705 82.915 89.875 83.085 ;
        RECT 90.165 82.915 90.335 83.085 ;
        RECT 90.625 82.915 90.795 83.085 ;
        RECT 91.085 82.915 91.255 83.085 ;
        RECT 91.545 82.915 91.715 83.085 ;
        RECT 92.005 82.915 92.175 83.085 ;
        RECT 92.465 82.915 92.635 83.085 ;
        RECT 92.925 82.915 93.095 83.085 ;
        RECT 93.385 82.915 93.555 83.085 ;
        RECT 93.845 82.915 94.015 83.085 ;
        RECT 94.305 82.915 94.475 83.085 ;
        RECT 94.765 82.915 94.935 83.085 ;
        RECT 95.225 82.915 95.395 83.085 ;
        RECT 95.685 82.915 95.855 83.085 ;
        RECT 96.145 82.915 96.315 83.085 ;
        RECT 96.605 82.915 96.775 83.085 ;
        RECT 97.065 82.915 97.235 83.085 ;
        RECT 97.525 82.915 97.695 83.085 ;
        RECT 97.985 82.915 98.155 83.085 ;
        RECT 98.445 82.915 98.615 83.085 ;
        RECT 98.905 82.915 99.075 83.085 ;
        RECT 99.365 82.915 99.535 83.085 ;
        RECT 99.825 82.915 99.995 83.085 ;
        RECT 100.285 82.915 100.455 83.085 ;
        RECT 100.745 82.915 100.915 83.085 ;
        RECT 101.205 82.915 101.375 83.085 ;
        RECT 101.665 82.915 101.835 83.085 ;
        RECT 102.125 82.915 102.295 83.085 ;
        RECT 102.585 82.915 102.755 83.085 ;
        RECT 103.045 82.915 103.215 83.085 ;
        RECT 103.505 82.915 103.675 83.085 ;
        RECT 103.965 82.915 104.135 83.085 ;
        RECT 104.425 82.915 104.595 83.085 ;
        RECT 104.885 82.915 105.055 83.085 ;
        RECT 105.345 82.915 105.515 83.085 ;
        RECT 105.805 82.915 105.975 83.085 ;
        RECT 106.265 82.915 106.435 83.085 ;
        RECT 106.725 82.915 106.895 83.085 ;
        RECT 107.185 82.915 107.355 83.085 ;
        RECT 107.645 82.915 107.815 83.085 ;
        RECT 108.105 82.915 108.275 83.085 ;
        RECT 108.565 82.915 108.735 83.085 ;
        RECT 109.025 82.915 109.195 83.085 ;
        RECT 109.485 82.915 109.655 83.085 ;
        RECT 109.945 82.915 110.115 83.085 ;
        RECT 110.405 82.915 110.575 83.085 ;
        RECT 110.865 82.915 111.035 83.085 ;
        RECT 111.325 82.915 111.495 83.085 ;
        RECT 111.785 82.915 111.955 83.085 ;
        RECT 112.245 82.915 112.415 83.085 ;
        RECT 112.705 82.915 112.875 83.085 ;
        RECT 113.165 82.915 113.335 83.085 ;
        RECT 113.625 82.915 113.795 83.085 ;
        RECT 114.085 82.915 114.255 83.085 ;
        RECT 114.545 82.915 114.715 83.085 ;
        RECT 115.005 82.915 115.175 83.085 ;
        RECT 115.465 82.915 115.635 83.085 ;
        RECT 115.925 82.915 116.095 83.085 ;
        RECT 116.385 82.915 116.555 83.085 ;
        RECT 116.845 82.915 117.015 83.085 ;
        RECT 117.305 82.915 117.475 83.085 ;
        RECT 117.765 82.915 117.935 83.085 ;
        RECT 118.225 82.915 118.395 83.085 ;
        RECT 118.685 82.915 118.855 83.085 ;
        RECT 119.145 82.915 119.315 83.085 ;
        RECT 119.605 82.915 119.775 83.085 ;
        RECT 120.065 82.915 120.235 83.085 ;
        RECT 120.525 82.915 120.695 83.085 ;
        RECT 120.985 82.915 121.155 83.085 ;
        RECT 121.445 82.915 121.615 83.085 ;
        RECT 121.905 82.915 122.075 83.085 ;
        RECT 122.365 82.915 122.535 83.085 ;
        RECT 122.825 82.915 122.995 83.085 ;
        RECT 123.285 82.915 123.455 83.085 ;
        RECT 123.745 82.915 123.915 83.085 ;
        RECT 124.205 82.915 124.375 83.085 ;
        RECT 124.665 82.915 124.835 83.085 ;
        RECT 125.125 82.915 125.295 83.085 ;
        RECT 125.585 82.915 125.755 83.085 ;
        RECT 126.045 82.915 126.215 83.085 ;
        RECT 126.505 82.915 126.675 83.085 ;
        RECT 126.965 82.915 127.135 83.085 ;
        RECT 127.425 82.915 127.595 83.085 ;
        RECT 127.885 82.915 128.055 83.085 ;
        RECT 128.345 82.915 128.515 83.085 ;
        RECT 128.805 82.915 128.975 83.085 ;
        RECT 129.265 82.915 129.435 83.085 ;
        RECT 129.725 82.915 129.895 83.085 ;
        RECT 130.185 82.915 130.355 83.085 ;
        RECT 130.645 82.915 130.815 83.085 ;
        RECT 131.105 82.915 131.275 83.085 ;
        RECT 131.565 82.915 131.735 83.085 ;
        RECT 132.025 82.915 132.195 83.085 ;
        RECT 132.485 82.915 132.655 83.085 ;
        RECT 132.945 82.915 133.115 83.085 ;
        RECT 133.405 82.915 133.575 83.085 ;
        RECT 133.865 82.915 134.035 83.085 ;
        RECT 134.325 82.915 134.495 83.085 ;
        RECT 134.785 82.915 134.955 83.085 ;
        RECT 135.245 82.915 135.415 83.085 ;
        RECT 135.705 82.915 135.875 83.085 ;
        RECT 136.165 82.915 136.335 83.085 ;
        RECT 136.625 82.915 136.795 83.085 ;
        RECT 137.085 82.915 137.255 83.085 ;
        RECT 137.545 82.915 137.715 83.085 ;
        RECT 138.005 82.915 138.175 83.085 ;
        RECT 138.465 82.915 138.635 83.085 ;
        RECT 138.925 82.915 139.095 83.085 ;
        RECT 139.385 82.915 139.555 83.085 ;
        RECT 139.845 82.915 140.015 83.085 ;
        RECT 140.305 82.915 140.475 83.085 ;
        RECT 140.765 82.915 140.935 83.085 ;
        RECT 141.225 82.915 141.395 83.085 ;
        RECT 141.685 82.915 141.855 83.085 ;
        RECT 142.145 82.915 142.315 83.085 ;
        RECT 142.605 82.915 142.775 83.085 ;
        RECT 143.065 82.915 143.235 83.085 ;
        RECT 143.525 82.915 143.695 83.085 ;
        RECT 143.985 82.915 144.155 83.085 ;
        RECT 55.665 77.475 55.835 77.645 ;
        RECT 56.125 77.475 56.295 77.645 ;
        RECT 56.585 77.475 56.755 77.645 ;
        RECT 57.045 77.475 57.215 77.645 ;
        RECT 57.505 77.475 57.675 77.645 ;
        RECT 57.965 77.475 58.135 77.645 ;
        RECT 58.425 77.475 58.595 77.645 ;
        RECT 58.885 77.475 59.055 77.645 ;
        RECT 59.345 77.475 59.515 77.645 ;
        RECT 59.805 77.475 59.975 77.645 ;
        RECT 60.265 77.475 60.435 77.645 ;
        RECT 60.725 77.475 60.895 77.645 ;
        RECT 61.185 77.475 61.355 77.645 ;
        RECT 61.645 77.475 61.815 77.645 ;
        RECT 62.105 77.475 62.275 77.645 ;
        RECT 62.565 77.475 62.735 77.645 ;
        RECT 63.025 77.475 63.195 77.645 ;
        RECT 63.485 77.475 63.655 77.645 ;
        RECT 63.945 77.475 64.115 77.645 ;
        RECT 64.405 77.475 64.575 77.645 ;
        RECT 64.865 77.475 65.035 77.645 ;
        RECT 65.325 77.475 65.495 77.645 ;
        RECT 65.785 77.475 65.955 77.645 ;
        RECT 66.245 77.475 66.415 77.645 ;
        RECT 66.705 77.475 66.875 77.645 ;
        RECT 67.165 77.475 67.335 77.645 ;
        RECT 67.625 77.475 67.795 77.645 ;
        RECT 68.085 77.475 68.255 77.645 ;
        RECT 68.545 77.475 68.715 77.645 ;
        RECT 69.005 77.475 69.175 77.645 ;
        RECT 69.465 77.475 69.635 77.645 ;
        RECT 69.925 77.475 70.095 77.645 ;
        RECT 70.385 77.475 70.555 77.645 ;
        RECT 70.845 77.475 71.015 77.645 ;
        RECT 71.305 77.475 71.475 77.645 ;
        RECT 71.765 77.475 71.935 77.645 ;
        RECT 72.225 77.475 72.395 77.645 ;
        RECT 72.685 77.475 72.855 77.645 ;
        RECT 73.145 77.475 73.315 77.645 ;
        RECT 73.605 77.475 73.775 77.645 ;
        RECT 74.065 77.475 74.235 77.645 ;
        RECT 74.525 77.475 74.695 77.645 ;
        RECT 74.985 77.475 75.155 77.645 ;
        RECT 75.445 77.475 75.615 77.645 ;
        RECT 75.905 77.475 76.075 77.645 ;
        RECT 76.365 77.475 76.535 77.645 ;
        RECT 76.825 77.475 76.995 77.645 ;
        RECT 77.285 77.475 77.455 77.645 ;
        RECT 77.745 77.475 77.915 77.645 ;
        RECT 78.205 77.475 78.375 77.645 ;
        RECT 78.665 77.475 78.835 77.645 ;
        RECT 79.125 77.475 79.295 77.645 ;
        RECT 79.585 77.475 79.755 77.645 ;
        RECT 80.045 77.475 80.215 77.645 ;
        RECT 80.505 77.475 80.675 77.645 ;
        RECT 80.965 77.475 81.135 77.645 ;
        RECT 81.425 77.475 81.595 77.645 ;
        RECT 81.885 77.475 82.055 77.645 ;
        RECT 82.345 77.475 82.515 77.645 ;
        RECT 82.805 77.475 82.975 77.645 ;
        RECT 83.265 77.475 83.435 77.645 ;
        RECT 83.725 77.475 83.895 77.645 ;
        RECT 84.185 77.475 84.355 77.645 ;
        RECT 84.645 77.475 84.815 77.645 ;
        RECT 85.105 77.475 85.275 77.645 ;
        RECT 85.565 77.475 85.735 77.645 ;
        RECT 86.025 77.475 86.195 77.645 ;
        RECT 86.485 77.475 86.655 77.645 ;
        RECT 86.945 77.475 87.115 77.645 ;
        RECT 87.405 77.475 87.575 77.645 ;
        RECT 87.865 77.475 88.035 77.645 ;
        RECT 88.325 77.475 88.495 77.645 ;
        RECT 88.785 77.475 88.955 77.645 ;
        RECT 89.245 77.475 89.415 77.645 ;
        RECT 89.705 77.475 89.875 77.645 ;
        RECT 90.165 77.475 90.335 77.645 ;
        RECT 90.625 77.475 90.795 77.645 ;
        RECT 91.085 77.475 91.255 77.645 ;
        RECT 91.545 77.475 91.715 77.645 ;
        RECT 92.005 77.475 92.175 77.645 ;
        RECT 92.465 77.475 92.635 77.645 ;
        RECT 92.925 77.475 93.095 77.645 ;
        RECT 93.385 77.475 93.555 77.645 ;
        RECT 93.845 77.475 94.015 77.645 ;
        RECT 94.305 77.475 94.475 77.645 ;
        RECT 94.765 77.475 94.935 77.645 ;
        RECT 95.225 77.475 95.395 77.645 ;
        RECT 95.685 77.475 95.855 77.645 ;
        RECT 96.145 77.475 96.315 77.645 ;
        RECT 96.605 77.475 96.775 77.645 ;
        RECT 97.065 77.475 97.235 77.645 ;
        RECT 97.525 77.475 97.695 77.645 ;
        RECT 97.985 77.475 98.155 77.645 ;
        RECT 98.445 77.475 98.615 77.645 ;
        RECT 98.905 77.475 99.075 77.645 ;
        RECT 99.365 77.475 99.535 77.645 ;
        RECT 99.825 77.475 99.995 77.645 ;
        RECT 100.285 77.475 100.455 77.645 ;
        RECT 100.745 77.475 100.915 77.645 ;
        RECT 101.205 77.475 101.375 77.645 ;
        RECT 101.665 77.475 101.835 77.645 ;
        RECT 102.125 77.475 102.295 77.645 ;
        RECT 102.585 77.475 102.755 77.645 ;
        RECT 103.045 77.475 103.215 77.645 ;
        RECT 103.505 77.475 103.675 77.645 ;
        RECT 103.965 77.475 104.135 77.645 ;
        RECT 104.425 77.475 104.595 77.645 ;
        RECT 104.885 77.475 105.055 77.645 ;
        RECT 105.345 77.475 105.515 77.645 ;
        RECT 105.805 77.475 105.975 77.645 ;
        RECT 106.265 77.475 106.435 77.645 ;
        RECT 106.725 77.475 106.895 77.645 ;
        RECT 107.185 77.475 107.355 77.645 ;
        RECT 107.645 77.475 107.815 77.645 ;
        RECT 108.105 77.475 108.275 77.645 ;
        RECT 108.565 77.475 108.735 77.645 ;
        RECT 109.025 77.475 109.195 77.645 ;
        RECT 109.485 77.475 109.655 77.645 ;
        RECT 109.945 77.475 110.115 77.645 ;
        RECT 110.405 77.475 110.575 77.645 ;
        RECT 110.865 77.475 111.035 77.645 ;
        RECT 111.325 77.475 111.495 77.645 ;
        RECT 111.785 77.475 111.955 77.645 ;
        RECT 112.245 77.475 112.415 77.645 ;
        RECT 112.705 77.475 112.875 77.645 ;
        RECT 113.165 77.475 113.335 77.645 ;
        RECT 113.625 77.475 113.795 77.645 ;
        RECT 114.085 77.475 114.255 77.645 ;
        RECT 114.545 77.475 114.715 77.645 ;
        RECT 115.005 77.475 115.175 77.645 ;
        RECT 115.465 77.475 115.635 77.645 ;
        RECT 115.925 77.475 116.095 77.645 ;
        RECT 116.385 77.475 116.555 77.645 ;
        RECT 116.845 77.475 117.015 77.645 ;
        RECT 117.305 77.475 117.475 77.645 ;
        RECT 117.765 77.475 117.935 77.645 ;
        RECT 118.225 77.475 118.395 77.645 ;
        RECT 118.685 77.475 118.855 77.645 ;
        RECT 119.145 77.475 119.315 77.645 ;
        RECT 119.605 77.475 119.775 77.645 ;
        RECT 120.065 77.475 120.235 77.645 ;
        RECT 120.525 77.475 120.695 77.645 ;
        RECT 120.985 77.475 121.155 77.645 ;
        RECT 121.445 77.475 121.615 77.645 ;
        RECT 121.905 77.475 122.075 77.645 ;
        RECT 122.365 77.475 122.535 77.645 ;
        RECT 122.825 77.475 122.995 77.645 ;
        RECT 123.285 77.475 123.455 77.645 ;
        RECT 123.745 77.475 123.915 77.645 ;
        RECT 124.205 77.475 124.375 77.645 ;
        RECT 124.665 77.475 124.835 77.645 ;
        RECT 125.125 77.475 125.295 77.645 ;
        RECT 125.585 77.475 125.755 77.645 ;
        RECT 126.045 77.475 126.215 77.645 ;
        RECT 126.505 77.475 126.675 77.645 ;
        RECT 126.965 77.475 127.135 77.645 ;
        RECT 127.425 77.475 127.595 77.645 ;
        RECT 127.885 77.475 128.055 77.645 ;
        RECT 128.345 77.475 128.515 77.645 ;
        RECT 128.805 77.475 128.975 77.645 ;
        RECT 129.265 77.475 129.435 77.645 ;
        RECT 129.725 77.475 129.895 77.645 ;
        RECT 130.185 77.475 130.355 77.645 ;
        RECT 130.645 77.475 130.815 77.645 ;
        RECT 131.105 77.475 131.275 77.645 ;
        RECT 131.565 77.475 131.735 77.645 ;
        RECT 132.025 77.475 132.195 77.645 ;
        RECT 132.485 77.475 132.655 77.645 ;
        RECT 132.945 77.475 133.115 77.645 ;
        RECT 133.405 77.475 133.575 77.645 ;
        RECT 133.865 77.475 134.035 77.645 ;
        RECT 134.325 77.475 134.495 77.645 ;
        RECT 134.785 77.475 134.955 77.645 ;
        RECT 135.245 77.475 135.415 77.645 ;
        RECT 135.705 77.475 135.875 77.645 ;
        RECT 136.165 77.475 136.335 77.645 ;
        RECT 136.625 77.475 136.795 77.645 ;
        RECT 137.085 77.475 137.255 77.645 ;
        RECT 137.545 77.475 137.715 77.645 ;
        RECT 138.005 77.475 138.175 77.645 ;
        RECT 138.465 77.475 138.635 77.645 ;
        RECT 138.925 77.475 139.095 77.645 ;
        RECT 139.385 77.475 139.555 77.645 ;
        RECT 139.845 77.475 140.015 77.645 ;
        RECT 140.305 77.475 140.475 77.645 ;
        RECT 140.765 77.475 140.935 77.645 ;
        RECT 141.225 77.475 141.395 77.645 ;
        RECT 141.685 77.475 141.855 77.645 ;
        RECT 142.145 77.475 142.315 77.645 ;
        RECT 142.605 77.475 142.775 77.645 ;
        RECT 143.065 77.475 143.235 77.645 ;
        RECT 143.525 77.475 143.695 77.645 ;
        RECT 143.985 77.475 144.155 77.645 ;
        RECT 55.665 72.035 55.835 72.205 ;
        RECT 56.125 72.035 56.295 72.205 ;
        RECT 56.585 72.035 56.755 72.205 ;
        RECT 57.045 72.035 57.215 72.205 ;
        RECT 57.505 72.035 57.675 72.205 ;
        RECT 57.965 72.035 58.135 72.205 ;
        RECT 58.425 72.035 58.595 72.205 ;
        RECT 58.885 72.035 59.055 72.205 ;
        RECT 59.345 72.035 59.515 72.205 ;
        RECT 59.805 72.035 59.975 72.205 ;
        RECT 60.265 72.035 60.435 72.205 ;
        RECT 60.725 72.035 60.895 72.205 ;
        RECT 61.185 72.035 61.355 72.205 ;
        RECT 61.645 72.035 61.815 72.205 ;
        RECT 62.105 72.035 62.275 72.205 ;
        RECT 62.565 72.035 62.735 72.205 ;
        RECT 63.025 72.035 63.195 72.205 ;
        RECT 63.485 72.035 63.655 72.205 ;
        RECT 63.945 72.035 64.115 72.205 ;
        RECT 64.405 72.035 64.575 72.205 ;
        RECT 64.865 72.035 65.035 72.205 ;
        RECT 65.325 72.035 65.495 72.205 ;
        RECT 65.785 72.035 65.955 72.205 ;
        RECT 66.245 72.035 66.415 72.205 ;
        RECT 66.705 72.035 66.875 72.205 ;
        RECT 67.165 72.035 67.335 72.205 ;
        RECT 67.625 72.035 67.795 72.205 ;
        RECT 68.085 72.035 68.255 72.205 ;
        RECT 68.545 72.035 68.715 72.205 ;
        RECT 69.005 72.035 69.175 72.205 ;
        RECT 69.465 72.035 69.635 72.205 ;
        RECT 69.925 72.035 70.095 72.205 ;
        RECT 70.385 72.035 70.555 72.205 ;
        RECT 70.845 72.035 71.015 72.205 ;
        RECT 71.305 72.035 71.475 72.205 ;
        RECT 71.765 72.035 71.935 72.205 ;
        RECT 72.225 72.035 72.395 72.205 ;
        RECT 72.685 72.035 72.855 72.205 ;
        RECT 73.145 72.035 73.315 72.205 ;
        RECT 73.605 72.035 73.775 72.205 ;
        RECT 74.065 72.035 74.235 72.205 ;
        RECT 74.525 72.035 74.695 72.205 ;
        RECT 74.985 72.035 75.155 72.205 ;
        RECT 75.445 72.035 75.615 72.205 ;
        RECT 75.905 72.035 76.075 72.205 ;
        RECT 76.365 72.035 76.535 72.205 ;
        RECT 76.825 72.035 76.995 72.205 ;
        RECT 77.285 72.035 77.455 72.205 ;
        RECT 77.745 72.035 77.915 72.205 ;
        RECT 78.205 72.035 78.375 72.205 ;
        RECT 78.665 72.035 78.835 72.205 ;
        RECT 79.125 72.035 79.295 72.205 ;
        RECT 79.585 72.035 79.755 72.205 ;
        RECT 80.045 72.035 80.215 72.205 ;
        RECT 80.505 72.035 80.675 72.205 ;
        RECT 80.965 72.035 81.135 72.205 ;
        RECT 81.425 72.035 81.595 72.205 ;
        RECT 81.885 72.035 82.055 72.205 ;
        RECT 82.345 72.035 82.515 72.205 ;
        RECT 82.805 72.035 82.975 72.205 ;
        RECT 83.265 72.035 83.435 72.205 ;
        RECT 83.725 72.035 83.895 72.205 ;
        RECT 84.185 72.035 84.355 72.205 ;
        RECT 84.645 72.035 84.815 72.205 ;
        RECT 85.105 72.035 85.275 72.205 ;
        RECT 85.565 72.035 85.735 72.205 ;
        RECT 86.025 72.035 86.195 72.205 ;
        RECT 86.485 72.035 86.655 72.205 ;
        RECT 86.945 72.035 87.115 72.205 ;
        RECT 87.405 72.035 87.575 72.205 ;
        RECT 87.865 72.035 88.035 72.205 ;
        RECT 88.325 72.035 88.495 72.205 ;
        RECT 88.785 72.035 88.955 72.205 ;
        RECT 89.245 72.035 89.415 72.205 ;
        RECT 89.705 72.035 89.875 72.205 ;
        RECT 90.165 72.035 90.335 72.205 ;
        RECT 90.625 72.035 90.795 72.205 ;
        RECT 91.085 72.035 91.255 72.205 ;
        RECT 91.545 72.035 91.715 72.205 ;
        RECT 92.005 72.035 92.175 72.205 ;
        RECT 92.465 72.035 92.635 72.205 ;
        RECT 92.925 72.035 93.095 72.205 ;
        RECT 93.385 72.035 93.555 72.205 ;
        RECT 93.845 72.035 94.015 72.205 ;
        RECT 94.305 72.035 94.475 72.205 ;
        RECT 94.765 72.035 94.935 72.205 ;
        RECT 95.225 72.035 95.395 72.205 ;
        RECT 95.685 72.035 95.855 72.205 ;
        RECT 96.145 72.035 96.315 72.205 ;
        RECT 96.605 72.035 96.775 72.205 ;
        RECT 97.065 72.035 97.235 72.205 ;
        RECT 97.525 72.035 97.695 72.205 ;
        RECT 97.985 72.035 98.155 72.205 ;
        RECT 98.445 72.035 98.615 72.205 ;
        RECT 98.905 72.035 99.075 72.205 ;
        RECT 99.365 72.035 99.535 72.205 ;
        RECT 99.825 72.035 99.995 72.205 ;
        RECT 100.285 72.035 100.455 72.205 ;
        RECT 100.745 72.035 100.915 72.205 ;
        RECT 101.205 72.035 101.375 72.205 ;
        RECT 101.665 72.035 101.835 72.205 ;
        RECT 102.125 72.035 102.295 72.205 ;
        RECT 102.585 72.035 102.755 72.205 ;
        RECT 103.045 72.035 103.215 72.205 ;
        RECT 103.505 72.035 103.675 72.205 ;
        RECT 103.965 72.035 104.135 72.205 ;
        RECT 104.425 72.035 104.595 72.205 ;
        RECT 104.885 72.035 105.055 72.205 ;
        RECT 105.345 72.035 105.515 72.205 ;
        RECT 105.805 72.035 105.975 72.205 ;
        RECT 106.265 72.035 106.435 72.205 ;
        RECT 106.725 72.035 106.895 72.205 ;
        RECT 107.185 72.035 107.355 72.205 ;
        RECT 107.645 72.035 107.815 72.205 ;
        RECT 108.105 72.035 108.275 72.205 ;
        RECT 108.565 72.035 108.735 72.205 ;
        RECT 109.025 72.035 109.195 72.205 ;
        RECT 109.485 72.035 109.655 72.205 ;
        RECT 109.945 72.035 110.115 72.205 ;
        RECT 110.405 72.035 110.575 72.205 ;
        RECT 110.865 72.035 111.035 72.205 ;
        RECT 111.325 72.035 111.495 72.205 ;
        RECT 111.785 72.035 111.955 72.205 ;
        RECT 112.245 72.035 112.415 72.205 ;
        RECT 112.705 72.035 112.875 72.205 ;
        RECT 113.165 72.035 113.335 72.205 ;
        RECT 113.625 72.035 113.795 72.205 ;
        RECT 114.085 72.035 114.255 72.205 ;
        RECT 114.545 72.035 114.715 72.205 ;
        RECT 115.005 72.035 115.175 72.205 ;
        RECT 115.465 72.035 115.635 72.205 ;
        RECT 115.925 72.035 116.095 72.205 ;
        RECT 116.385 72.035 116.555 72.205 ;
        RECT 116.845 72.035 117.015 72.205 ;
        RECT 117.305 72.035 117.475 72.205 ;
        RECT 117.765 72.035 117.935 72.205 ;
        RECT 118.225 72.035 118.395 72.205 ;
        RECT 118.685 72.035 118.855 72.205 ;
        RECT 119.145 72.035 119.315 72.205 ;
        RECT 119.605 72.035 119.775 72.205 ;
        RECT 120.065 72.035 120.235 72.205 ;
        RECT 120.525 72.035 120.695 72.205 ;
        RECT 120.985 72.035 121.155 72.205 ;
        RECT 121.445 72.035 121.615 72.205 ;
        RECT 121.905 72.035 122.075 72.205 ;
        RECT 122.365 72.035 122.535 72.205 ;
        RECT 122.825 72.035 122.995 72.205 ;
        RECT 123.285 72.035 123.455 72.205 ;
        RECT 123.745 72.035 123.915 72.205 ;
        RECT 124.205 72.035 124.375 72.205 ;
        RECT 124.665 72.035 124.835 72.205 ;
        RECT 125.125 72.035 125.295 72.205 ;
        RECT 125.585 72.035 125.755 72.205 ;
        RECT 126.045 72.035 126.215 72.205 ;
        RECT 126.505 72.035 126.675 72.205 ;
        RECT 126.965 72.035 127.135 72.205 ;
        RECT 127.425 72.035 127.595 72.205 ;
        RECT 127.885 72.035 128.055 72.205 ;
        RECT 128.345 72.035 128.515 72.205 ;
        RECT 128.805 72.035 128.975 72.205 ;
        RECT 129.265 72.035 129.435 72.205 ;
        RECT 129.725 72.035 129.895 72.205 ;
        RECT 130.185 72.035 130.355 72.205 ;
        RECT 130.645 72.035 130.815 72.205 ;
        RECT 131.105 72.035 131.275 72.205 ;
        RECT 131.565 72.035 131.735 72.205 ;
        RECT 132.025 72.035 132.195 72.205 ;
        RECT 132.485 72.035 132.655 72.205 ;
        RECT 132.945 72.035 133.115 72.205 ;
        RECT 133.405 72.035 133.575 72.205 ;
        RECT 133.865 72.035 134.035 72.205 ;
        RECT 134.325 72.035 134.495 72.205 ;
        RECT 134.785 72.035 134.955 72.205 ;
        RECT 135.245 72.035 135.415 72.205 ;
        RECT 135.705 72.035 135.875 72.205 ;
        RECT 136.165 72.035 136.335 72.205 ;
        RECT 136.625 72.035 136.795 72.205 ;
        RECT 137.085 72.035 137.255 72.205 ;
        RECT 137.545 72.035 137.715 72.205 ;
        RECT 138.005 72.035 138.175 72.205 ;
        RECT 138.465 72.035 138.635 72.205 ;
        RECT 138.925 72.035 139.095 72.205 ;
        RECT 139.385 72.035 139.555 72.205 ;
        RECT 139.845 72.035 140.015 72.205 ;
        RECT 140.305 72.035 140.475 72.205 ;
        RECT 140.765 72.035 140.935 72.205 ;
        RECT 141.225 72.035 141.395 72.205 ;
        RECT 141.685 72.035 141.855 72.205 ;
        RECT 142.145 72.035 142.315 72.205 ;
        RECT 142.605 72.035 142.775 72.205 ;
        RECT 143.065 72.035 143.235 72.205 ;
        RECT 143.525 72.035 143.695 72.205 ;
        RECT 143.985 72.035 144.155 72.205 ;
        RECT 55.665 66.595 55.835 66.765 ;
        RECT 56.125 66.595 56.295 66.765 ;
        RECT 56.585 66.595 56.755 66.765 ;
        RECT 57.045 66.595 57.215 66.765 ;
        RECT 57.505 66.595 57.675 66.765 ;
        RECT 57.965 66.595 58.135 66.765 ;
        RECT 58.425 66.595 58.595 66.765 ;
        RECT 58.885 66.595 59.055 66.765 ;
        RECT 59.345 66.595 59.515 66.765 ;
        RECT 59.805 66.595 59.975 66.765 ;
        RECT 60.265 66.595 60.435 66.765 ;
        RECT 60.725 66.595 60.895 66.765 ;
        RECT 61.185 66.595 61.355 66.765 ;
        RECT 61.645 66.595 61.815 66.765 ;
        RECT 62.105 66.595 62.275 66.765 ;
        RECT 62.565 66.595 62.735 66.765 ;
        RECT 63.025 66.595 63.195 66.765 ;
        RECT 63.485 66.595 63.655 66.765 ;
        RECT 63.945 66.595 64.115 66.765 ;
        RECT 64.405 66.595 64.575 66.765 ;
        RECT 64.865 66.595 65.035 66.765 ;
        RECT 65.325 66.595 65.495 66.765 ;
        RECT 65.785 66.595 65.955 66.765 ;
        RECT 66.245 66.595 66.415 66.765 ;
        RECT 66.705 66.595 66.875 66.765 ;
        RECT 67.165 66.595 67.335 66.765 ;
        RECT 67.625 66.595 67.795 66.765 ;
        RECT 68.085 66.595 68.255 66.765 ;
        RECT 68.545 66.595 68.715 66.765 ;
        RECT 69.005 66.595 69.175 66.765 ;
        RECT 69.465 66.595 69.635 66.765 ;
        RECT 69.925 66.595 70.095 66.765 ;
        RECT 70.385 66.595 70.555 66.765 ;
        RECT 70.845 66.595 71.015 66.765 ;
        RECT 71.305 66.595 71.475 66.765 ;
        RECT 71.765 66.595 71.935 66.765 ;
        RECT 72.225 66.595 72.395 66.765 ;
        RECT 72.685 66.595 72.855 66.765 ;
        RECT 73.145 66.595 73.315 66.765 ;
        RECT 73.605 66.595 73.775 66.765 ;
        RECT 74.065 66.595 74.235 66.765 ;
        RECT 74.525 66.595 74.695 66.765 ;
        RECT 74.985 66.595 75.155 66.765 ;
        RECT 75.445 66.595 75.615 66.765 ;
        RECT 75.905 66.595 76.075 66.765 ;
        RECT 76.365 66.595 76.535 66.765 ;
        RECT 76.825 66.595 76.995 66.765 ;
        RECT 77.285 66.595 77.455 66.765 ;
        RECT 77.745 66.595 77.915 66.765 ;
        RECT 78.205 66.595 78.375 66.765 ;
        RECT 78.665 66.595 78.835 66.765 ;
        RECT 79.125 66.595 79.295 66.765 ;
        RECT 79.585 66.595 79.755 66.765 ;
        RECT 80.045 66.595 80.215 66.765 ;
        RECT 80.505 66.595 80.675 66.765 ;
        RECT 80.965 66.595 81.135 66.765 ;
        RECT 81.425 66.595 81.595 66.765 ;
        RECT 81.885 66.595 82.055 66.765 ;
        RECT 82.345 66.595 82.515 66.765 ;
        RECT 82.805 66.595 82.975 66.765 ;
        RECT 83.265 66.595 83.435 66.765 ;
        RECT 83.725 66.595 83.895 66.765 ;
        RECT 84.185 66.595 84.355 66.765 ;
        RECT 84.645 66.595 84.815 66.765 ;
        RECT 85.105 66.595 85.275 66.765 ;
        RECT 85.565 66.595 85.735 66.765 ;
        RECT 86.025 66.595 86.195 66.765 ;
        RECT 86.485 66.595 86.655 66.765 ;
        RECT 86.945 66.595 87.115 66.765 ;
        RECT 87.405 66.595 87.575 66.765 ;
        RECT 87.865 66.595 88.035 66.765 ;
        RECT 88.325 66.595 88.495 66.765 ;
        RECT 88.785 66.595 88.955 66.765 ;
        RECT 89.245 66.595 89.415 66.765 ;
        RECT 89.705 66.595 89.875 66.765 ;
        RECT 90.165 66.595 90.335 66.765 ;
        RECT 90.625 66.595 90.795 66.765 ;
        RECT 91.085 66.595 91.255 66.765 ;
        RECT 91.545 66.595 91.715 66.765 ;
        RECT 92.005 66.595 92.175 66.765 ;
        RECT 92.465 66.595 92.635 66.765 ;
        RECT 92.925 66.595 93.095 66.765 ;
        RECT 93.385 66.595 93.555 66.765 ;
        RECT 93.845 66.595 94.015 66.765 ;
        RECT 94.305 66.595 94.475 66.765 ;
        RECT 94.765 66.595 94.935 66.765 ;
        RECT 95.225 66.595 95.395 66.765 ;
        RECT 95.685 66.595 95.855 66.765 ;
        RECT 96.145 66.595 96.315 66.765 ;
        RECT 96.605 66.595 96.775 66.765 ;
        RECT 97.065 66.595 97.235 66.765 ;
        RECT 97.525 66.595 97.695 66.765 ;
        RECT 97.985 66.595 98.155 66.765 ;
        RECT 98.445 66.595 98.615 66.765 ;
        RECT 98.905 66.595 99.075 66.765 ;
        RECT 99.365 66.595 99.535 66.765 ;
        RECT 99.825 66.595 99.995 66.765 ;
        RECT 100.285 66.595 100.455 66.765 ;
        RECT 100.745 66.595 100.915 66.765 ;
        RECT 101.205 66.595 101.375 66.765 ;
        RECT 101.665 66.595 101.835 66.765 ;
        RECT 102.125 66.595 102.295 66.765 ;
        RECT 102.585 66.595 102.755 66.765 ;
        RECT 103.045 66.595 103.215 66.765 ;
        RECT 103.505 66.595 103.675 66.765 ;
        RECT 103.965 66.595 104.135 66.765 ;
        RECT 104.425 66.595 104.595 66.765 ;
        RECT 104.885 66.595 105.055 66.765 ;
        RECT 105.345 66.595 105.515 66.765 ;
        RECT 105.805 66.595 105.975 66.765 ;
        RECT 106.265 66.595 106.435 66.765 ;
        RECT 106.725 66.595 106.895 66.765 ;
        RECT 107.185 66.595 107.355 66.765 ;
        RECT 107.645 66.595 107.815 66.765 ;
        RECT 108.105 66.595 108.275 66.765 ;
        RECT 108.565 66.595 108.735 66.765 ;
        RECT 109.025 66.595 109.195 66.765 ;
        RECT 109.485 66.595 109.655 66.765 ;
        RECT 109.945 66.595 110.115 66.765 ;
        RECT 110.405 66.595 110.575 66.765 ;
        RECT 110.865 66.595 111.035 66.765 ;
        RECT 111.325 66.595 111.495 66.765 ;
        RECT 111.785 66.595 111.955 66.765 ;
        RECT 112.245 66.595 112.415 66.765 ;
        RECT 112.705 66.595 112.875 66.765 ;
        RECT 113.165 66.595 113.335 66.765 ;
        RECT 113.625 66.595 113.795 66.765 ;
        RECT 114.085 66.595 114.255 66.765 ;
        RECT 114.545 66.595 114.715 66.765 ;
        RECT 115.005 66.595 115.175 66.765 ;
        RECT 115.465 66.595 115.635 66.765 ;
        RECT 115.925 66.595 116.095 66.765 ;
        RECT 116.385 66.595 116.555 66.765 ;
        RECT 116.845 66.595 117.015 66.765 ;
        RECT 117.305 66.595 117.475 66.765 ;
        RECT 117.765 66.595 117.935 66.765 ;
        RECT 118.225 66.595 118.395 66.765 ;
        RECT 118.685 66.595 118.855 66.765 ;
        RECT 119.145 66.595 119.315 66.765 ;
        RECT 119.605 66.595 119.775 66.765 ;
        RECT 120.065 66.595 120.235 66.765 ;
        RECT 120.525 66.595 120.695 66.765 ;
        RECT 120.985 66.595 121.155 66.765 ;
        RECT 121.445 66.595 121.615 66.765 ;
        RECT 121.905 66.595 122.075 66.765 ;
        RECT 122.365 66.595 122.535 66.765 ;
        RECT 122.825 66.595 122.995 66.765 ;
        RECT 123.285 66.595 123.455 66.765 ;
        RECT 123.745 66.595 123.915 66.765 ;
        RECT 124.205 66.595 124.375 66.765 ;
        RECT 124.665 66.595 124.835 66.765 ;
        RECT 125.125 66.595 125.295 66.765 ;
        RECT 125.585 66.595 125.755 66.765 ;
        RECT 126.045 66.595 126.215 66.765 ;
        RECT 126.505 66.595 126.675 66.765 ;
        RECT 126.965 66.595 127.135 66.765 ;
        RECT 127.425 66.595 127.595 66.765 ;
        RECT 127.885 66.595 128.055 66.765 ;
        RECT 128.345 66.595 128.515 66.765 ;
        RECT 128.805 66.595 128.975 66.765 ;
        RECT 129.265 66.595 129.435 66.765 ;
        RECT 129.725 66.595 129.895 66.765 ;
        RECT 130.185 66.595 130.355 66.765 ;
        RECT 130.645 66.595 130.815 66.765 ;
        RECT 131.105 66.595 131.275 66.765 ;
        RECT 131.565 66.595 131.735 66.765 ;
        RECT 132.025 66.595 132.195 66.765 ;
        RECT 132.485 66.595 132.655 66.765 ;
        RECT 132.945 66.595 133.115 66.765 ;
        RECT 133.405 66.595 133.575 66.765 ;
        RECT 133.865 66.595 134.035 66.765 ;
        RECT 134.325 66.595 134.495 66.765 ;
        RECT 134.785 66.595 134.955 66.765 ;
        RECT 135.245 66.595 135.415 66.765 ;
        RECT 135.705 66.595 135.875 66.765 ;
        RECT 136.165 66.595 136.335 66.765 ;
        RECT 136.625 66.595 136.795 66.765 ;
        RECT 137.085 66.595 137.255 66.765 ;
        RECT 137.545 66.595 137.715 66.765 ;
        RECT 138.005 66.595 138.175 66.765 ;
        RECT 138.465 66.595 138.635 66.765 ;
        RECT 138.925 66.595 139.095 66.765 ;
        RECT 139.385 66.595 139.555 66.765 ;
        RECT 139.845 66.595 140.015 66.765 ;
        RECT 140.305 66.595 140.475 66.765 ;
        RECT 140.765 66.595 140.935 66.765 ;
        RECT 141.225 66.595 141.395 66.765 ;
        RECT 141.685 66.595 141.855 66.765 ;
        RECT 142.145 66.595 142.315 66.765 ;
        RECT 142.605 66.595 142.775 66.765 ;
        RECT 143.065 66.595 143.235 66.765 ;
        RECT 143.525 66.595 143.695 66.765 ;
        RECT 143.985 66.595 144.155 66.765 ;
        RECT 55.665 61.155 55.835 61.325 ;
        RECT 56.125 61.155 56.295 61.325 ;
        RECT 56.585 61.155 56.755 61.325 ;
        RECT 57.045 61.155 57.215 61.325 ;
        RECT 57.505 61.155 57.675 61.325 ;
        RECT 57.965 61.155 58.135 61.325 ;
        RECT 58.425 61.155 58.595 61.325 ;
        RECT 58.885 61.155 59.055 61.325 ;
        RECT 59.345 61.155 59.515 61.325 ;
        RECT 59.805 61.155 59.975 61.325 ;
        RECT 60.265 61.155 60.435 61.325 ;
        RECT 60.725 61.155 60.895 61.325 ;
        RECT 61.185 61.155 61.355 61.325 ;
        RECT 61.645 61.155 61.815 61.325 ;
        RECT 62.105 61.155 62.275 61.325 ;
        RECT 62.565 61.155 62.735 61.325 ;
        RECT 63.025 61.155 63.195 61.325 ;
        RECT 63.485 61.155 63.655 61.325 ;
        RECT 63.945 61.155 64.115 61.325 ;
        RECT 64.405 61.155 64.575 61.325 ;
        RECT 64.865 61.155 65.035 61.325 ;
        RECT 65.325 61.155 65.495 61.325 ;
        RECT 65.785 61.155 65.955 61.325 ;
        RECT 66.245 61.155 66.415 61.325 ;
        RECT 66.705 61.155 66.875 61.325 ;
        RECT 67.165 61.155 67.335 61.325 ;
        RECT 67.625 61.155 67.795 61.325 ;
        RECT 68.085 61.155 68.255 61.325 ;
        RECT 68.545 61.155 68.715 61.325 ;
        RECT 69.005 61.155 69.175 61.325 ;
        RECT 69.465 61.155 69.635 61.325 ;
        RECT 69.925 61.155 70.095 61.325 ;
        RECT 70.385 61.155 70.555 61.325 ;
        RECT 70.845 61.155 71.015 61.325 ;
        RECT 71.305 61.155 71.475 61.325 ;
        RECT 71.765 61.155 71.935 61.325 ;
        RECT 72.225 61.155 72.395 61.325 ;
        RECT 72.685 61.155 72.855 61.325 ;
        RECT 73.145 61.155 73.315 61.325 ;
        RECT 73.605 61.155 73.775 61.325 ;
        RECT 74.065 61.155 74.235 61.325 ;
        RECT 74.525 61.155 74.695 61.325 ;
        RECT 74.985 61.155 75.155 61.325 ;
        RECT 75.445 61.155 75.615 61.325 ;
        RECT 75.905 61.155 76.075 61.325 ;
        RECT 76.365 61.155 76.535 61.325 ;
        RECT 76.825 61.155 76.995 61.325 ;
        RECT 77.285 61.155 77.455 61.325 ;
        RECT 77.745 61.155 77.915 61.325 ;
        RECT 78.205 61.155 78.375 61.325 ;
        RECT 78.665 61.155 78.835 61.325 ;
        RECT 79.125 61.155 79.295 61.325 ;
        RECT 79.585 61.155 79.755 61.325 ;
        RECT 80.045 61.155 80.215 61.325 ;
        RECT 80.505 61.155 80.675 61.325 ;
        RECT 80.965 61.155 81.135 61.325 ;
        RECT 81.425 61.155 81.595 61.325 ;
        RECT 81.885 61.155 82.055 61.325 ;
        RECT 82.345 61.155 82.515 61.325 ;
        RECT 82.805 61.155 82.975 61.325 ;
        RECT 83.265 61.155 83.435 61.325 ;
        RECT 83.725 61.155 83.895 61.325 ;
        RECT 84.185 61.155 84.355 61.325 ;
        RECT 84.645 61.155 84.815 61.325 ;
        RECT 85.105 61.155 85.275 61.325 ;
        RECT 85.565 61.155 85.735 61.325 ;
        RECT 86.025 61.155 86.195 61.325 ;
        RECT 86.485 61.155 86.655 61.325 ;
        RECT 86.945 61.155 87.115 61.325 ;
        RECT 87.405 61.155 87.575 61.325 ;
        RECT 87.865 61.155 88.035 61.325 ;
        RECT 88.325 61.155 88.495 61.325 ;
        RECT 88.785 61.155 88.955 61.325 ;
        RECT 89.245 61.155 89.415 61.325 ;
        RECT 89.705 61.155 89.875 61.325 ;
        RECT 90.165 61.155 90.335 61.325 ;
        RECT 90.625 61.155 90.795 61.325 ;
        RECT 91.085 61.155 91.255 61.325 ;
        RECT 91.545 61.155 91.715 61.325 ;
        RECT 92.005 61.155 92.175 61.325 ;
        RECT 92.465 61.155 92.635 61.325 ;
        RECT 92.925 61.155 93.095 61.325 ;
        RECT 93.385 61.155 93.555 61.325 ;
        RECT 93.845 61.155 94.015 61.325 ;
        RECT 94.305 61.155 94.475 61.325 ;
        RECT 94.765 61.155 94.935 61.325 ;
        RECT 95.225 61.155 95.395 61.325 ;
        RECT 95.685 61.155 95.855 61.325 ;
        RECT 96.145 61.155 96.315 61.325 ;
        RECT 96.605 61.155 96.775 61.325 ;
        RECT 97.065 61.155 97.235 61.325 ;
        RECT 97.525 61.155 97.695 61.325 ;
        RECT 97.985 61.155 98.155 61.325 ;
        RECT 98.445 61.155 98.615 61.325 ;
        RECT 98.905 61.155 99.075 61.325 ;
        RECT 99.365 61.155 99.535 61.325 ;
        RECT 99.825 61.155 99.995 61.325 ;
        RECT 100.285 61.155 100.455 61.325 ;
        RECT 100.745 61.155 100.915 61.325 ;
        RECT 101.205 61.155 101.375 61.325 ;
        RECT 101.665 61.155 101.835 61.325 ;
        RECT 102.125 61.155 102.295 61.325 ;
        RECT 102.585 61.155 102.755 61.325 ;
        RECT 103.045 61.155 103.215 61.325 ;
        RECT 103.505 61.155 103.675 61.325 ;
        RECT 103.965 61.155 104.135 61.325 ;
        RECT 104.425 61.155 104.595 61.325 ;
        RECT 104.885 61.155 105.055 61.325 ;
        RECT 105.345 61.155 105.515 61.325 ;
        RECT 105.805 61.155 105.975 61.325 ;
        RECT 106.265 61.155 106.435 61.325 ;
        RECT 106.725 61.155 106.895 61.325 ;
        RECT 107.185 61.155 107.355 61.325 ;
        RECT 107.645 61.155 107.815 61.325 ;
        RECT 108.105 61.155 108.275 61.325 ;
        RECT 108.565 61.155 108.735 61.325 ;
        RECT 109.025 61.155 109.195 61.325 ;
        RECT 109.485 61.155 109.655 61.325 ;
        RECT 109.945 61.155 110.115 61.325 ;
        RECT 110.405 61.155 110.575 61.325 ;
        RECT 110.865 61.155 111.035 61.325 ;
        RECT 111.325 61.155 111.495 61.325 ;
        RECT 111.785 61.155 111.955 61.325 ;
        RECT 112.245 61.155 112.415 61.325 ;
        RECT 112.705 61.155 112.875 61.325 ;
        RECT 113.165 61.155 113.335 61.325 ;
        RECT 113.625 61.155 113.795 61.325 ;
        RECT 114.085 61.155 114.255 61.325 ;
        RECT 114.545 61.155 114.715 61.325 ;
        RECT 115.005 61.155 115.175 61.325 ;
        RECT 115.465 61.155 115.635 61.325 ;
        RECT 115.925 61.155 116.095 61.325 ;
        RECT 116.385 61.155 116.555 61.325 ;
        RECT 116.845 61.155 117.015 61.325 ;
        RECT 117.305 61.155 117.475 61.325 ;
        RECT 117.765 61.155 117.935 61.325 ;
        RECT 118.225 61.155 118.395 61.325 ;
        RECT 118.685 61.155 118.855 61.325 ;
        RECT 119.145 61.155 119.315 61.325 ;
        RECT 119.605 61.155 119.775 61.325 ;
        RECT 120.065 61.155 120.235 61.325 ;
        RECT 120.525 61.155 120.695 61.325 ;
        RECT 120.985 61.155 121.155 61.325 ;
        RECT 121.445 61.155 121.615 61.325 ;
        RECT 121.905 61.155 122.075 61.325 ;
        RECT 122.365 61.155 122.535 61.325 ;
        RECT 122.825 61.155 122.995 61.325 ;
        RECT 123.285 61.155 123.455 61.325 ;
        RECT 123.745 61.155 123.915 61.325 ;
        RECT 124.205 61.155 124.375 61.325 ;
        RECT 124.665 61.155 124.835 61.325 ;
        RECT 125.125 61.155 125.295 61.325 ;
        RECT 125.585 61.155 125.755 61.325 ;
        RECT 126.045 61.155 126.215 61.325 ;
        RECT 126.505 61.155 126.675 61.325 ;
        RECT 126.965 61.155 127.135 61.325 ;
        RECT 127.425 61.155 127.595 61.325 ;
        RECT 127.885 61.155 128.055 61.325 ;
        RECT 128.345 61.155 128.515 61.325 ;
        RECT 128.805 61.155 128.975 61.325 ;
        RECT 129.265 61.155 129.435 61.325 ;
        RECT 129.725 61.155 129.895 61.325 ;
        RECT 130.185 61.155 130.355 61.325 ;
        RECT 130.645 61.155 130.815 61.325 ;
        RECT 131.105 61.155 131.275 61.325 ;
        RECT 131.565 61.155 131.735 61.325 ;
        RECT 132.025 61.155 132.195 61.325 ;
        RECT 132.485 61.155 132.655 61.325 ;
        RECT 132.945 61.155 133.115 61.325 ;
        RECT 133.405 61.155 133.575 61.325 ;
        RECT 133.865 61.155 134.035 61.325 ;
        RECT 134.325 61.155 134.495 61.325 ;
        RECT 134.785 61.155 134.955 61.325 ;
        RECT 135.245 61.155 135.415 61.325 ;
        RECT 135.705 61.155 135.875 61.325 ;
        RECT 136.165 61.155 136.335 61.325 ;
        RECT 136.625 61.155 136.795 61.325 ;
        RECT 137.085 61.155 137.255 61.325 ;
        RECT 137.545 61.155 137.715 61.325 ;
        RECT 138.005 61.155 138.175 61.325 ;
        RECT 138.465 61.155 138.635 61.325 ;
        RECT 138.925 61.155 139.095 61.325 ;
        RECT 139.385 61.155 139.555 61.325 ;
        RECT 139.845 61.155 140.015 61.325 ;
        RECT 140.305 61.155 140.475 61.325 ;
        RECT 140.765 61.155 140.935 61.325 ;
        RECT 141.225 61.155 141.395 61.325 ;
        RECT 141.685 61.155 141.855 61.325 ;
        RECT 142.145 61.155 142.315 61.325 ;
        RECT 142.605 61.155 142.775 61.325 ;
        RECT 143.065 61.155 143.235 61.325 ;
        RECT 143.525 61.155 143.695 61.325 ;
        RECT 143.985 61.155 144.155 61.325 ;
        RECT 55.665 55.715 55.835 55.885 ;
        RECT 56.125 55.715 56.295 55.885 ;
        RECT 56.585 55.715 56.755 55.885 ;
        RECT 57.045 55.715 57.215 55.885 ;
        RECT 57.505 55.715 57.675 55.885 ;
        RECT 57.965 55.715 58.135 55.885 ;
        RECT 58.425 55.715 58.595 55.885 ;
        RECT 58.885 55.715 59.055 55.885 ;
        RECT 59.345 55.715 59.515 55.885 ;
        RECT 59.805 55.715 59.975 55.885 ;
        RECT 60.265 55.715 60.435 55.885 ;
        RECT 60.725 55.715 60.895 55.885 ;
        RECT 61.185 55.715 61.355 55.885 ;
        RECT 61.645 55.715 61.815 55.885 ;
        RECT 62.105 55.715 62.275 55.885 ;
        RECT 62.565 55.715 62.735 55.885 ;
        RECT 63.025 55.715 63.195 55.885 ;
        RECT 63.485 55.715 63.655 55.885 ;
        RECT 63.945 55.715 64.115 55.885 ;
        RECT 64.405 55.715 64.575 55.885 ;
        RECT 64.865 55.715 65.035 55.885 ;
        RECT 65.325 55.715 65.495 55.885 ;
        RECT 65.785 55.715 65.955 55.885 ;
        RECT 66.245 55.715 66.415 55.885 ;
        RECT 66.705 55.715 66.875 55.885 ;
        RECT 67.165 55.715 67.335 55.885 ;
        RECT 67.625 55.715 67.795 55.885 ;
        RECT 68.085 55.715 68.255 55.885 ;
        RECT 68.545 55.715 68.715 55.885 ;
        RECT 69.005 55.715 69.175 55.885 ;
        RECT 69.465 55.715 69.635 55.885 ;
        RECT 69.925 55.715 70.095 55.885 ;
        RECT 70.385 55.715 70.555 55.885 ;
        RECT 70.845 55.715 71.015 55.885 ;
        RECT 71.305 55.715 71.475 55.885 ;
        RECT 71.765 55.715 71.935 55.885 ;
        RECT 72.225 55.715 72.395 55.885 ;
        RECT 72.685 55.715 72.855 55.885 ;
        RECT 73.145 55.715 73.315 55.885 ;
        RECT 73.605 55.715 73.775 55.885 ;
        RECT 74.065 55.715 74.235 55.885 ;
        RECT 74.525 55.715 74.695 55.885 ;
        RECT 74.985 55.715 75.155 55.885 ;
        RECT 75.445 55.715 75.615 55.885 ;
        RECT 75.905 55.715 76.075 55.885 ;
        RECT 76.365 55.715 76.535 55.885 ;
        RECT 76.825 55.715 76.995 55.885 ;
        RECT 77.285 55.715 77.455 55.885 ;
        RECT 77.745 55.715 77.915 55.885 ;
        RECT 78.205 55.715 78.375 55.885 ;
        RECT 78.665 55.715 78.835 55.885 ;
        RECT 79.125 55.715 79.295 55.885 ;
        RECT 79.585 55.715 79.755 55.885 ;
        RECT 80.045 55.715 80.215 55.885 ;
        RECT 80.505 55.715 80.675 55.885 ;
        RECT 80.965 55.715 81.135 55.885 ;
        RECT 81.425 55.715 81.595 55.885 ;
        RECT 81.885 55.715 82.055 55.885 ;
        RECT 82.345 55.715 82.515 55.885 ;
        RECT 82.805 55.715 82.975 55.885 ;
        RECT 83.265 55.715 83.435 55.885 ;
        RECT 83.725 55.715 83.895 55.885 ;
        RECT 84.185 55.715 84.355 55.885 ;
        RECT 84.645 55.715 84.815 55.885 ;
        RECT 85.105 55.715 85.275 55.885 ;
        RECT 85.565 55.715 85.735 55.885 ;
        RECT 86.025 55.715 86.195 55.885 ;
        RECT 86.485 55.715 86.655 55.885 ;
        RECT 86.945 55.715 87.115 55.885 ;
        RECT 87.405 55.715 87.575 55.885 ;
        RECT 87.865 55.715 88.035 55.885 ;
        RECT 88.325 55.715 88.495 55.885 ;
        RECT 88.785 55.715 88.955 55.885 ;
        RECT 89.245 55.715 89.415 55.885 ;
        RECT 89.705 55.715 89.875 55.885 ;
        RECT 90.165 55.715 90.335 55.885 ;
        RECT 90.625 55.715 90.795 55.885 ;
        RECT 91.085 55.715 91.255 55.885 ;
        RECT 91.545 55.715 91.715 55.885 ;
        RECT 92.005 55.715 92.175 55.885 ;
        RECT 92.465 55.715 92.635 55.885 ;
        RECT 92.925 55.715 93.095 55.885 ;
        RECT 93.385 55.715 93.555 55.885 ;
        RECT 93.845 55.715 94.015 55.885 ;
        RECT 94.305 55.715 94.475 55.885 ;
        RECT 94.765 55.715 94.935 55.885 ;
        RECT 95.225 55.715 95.395 55.885 ;
        RECT 95.685 55.715 95.855 55.885 ;
        RECT 96.145 55.715 96.315 55.885 ;
        RECT 96.605 55.715 96.775 55.885 ;
        RECT 97.065 55.715 97.235 55.885 ;
        RECT 97.525 55.715 97.695 55.885 ;
        RECT 97.985 55.715 98.155 55.885 ;
        RECT 98.445 55.715 98.615 55.885 ;
        RECT 98.905 55.715 99.075 55.885 ;
        RECT 99.365 55.715 99.535 55.885 ;
        RECT 99.825 55.715 99.995 55.885 ;
        RECT 100.285 55.715 100.455 55.885 ;
        RECT 100.745 55.715 100.915 55.885 ;
        RECT 101.205 55.715 101.375 55.885 ;
        RECT 101.665 55.715 101.835 55.885 ;
        RECT 102.125 55.715 102.295 55.885 ;
        RECT 102.585 55.715 102.755 55.885 ;
        RECT 103.045 55.715 103.215 55.885 ;
        RECT 103.505 55.715 103.675 55.885 ;
        RECT 103.965 55.715 104.135 55.885 ;
        RECT 104.425 55.715 104.595 55.885 ;
        RECT 104.885 55.715 105.055 55.885 ;
        RECT 105.345 55.715 105.515 55.885 ;
        RECT 105.805 55.715 105.975 55.885 ;
        RECT 106.265 55.715 106.435 55.885 ;
        RECT 106.725 55.715 106.895 55.885 ;
        RECT 107.185 55.715 107.355 55.885 ;
        RECT 107.645 55.715 107.815 55.885 ;
        RECT 108.105 55.715 108.275 55.885 ;
        RECT 108.565 55.715 108.735 55.885 ;
        RECT 109.025 55.715 109.195 55.885 ;
        RECT 109.485 55.715 109.655 55.885 ;
        RECT 109.945 55.715 110.115 55.885 ;
        RECT 110.405 55.715 110.575 55.885 ;
        RECT 110.865 55.715 111.035 55.885 ;
        RECT 111.325 55.715 111.495 55.885 ;
        RECT 111.785 55.715 111.955 55.885 ;
        RECT 112.245 55.715 112.415 55.885 ;
        RECT 112.705 55.715 112.875 55.885 ;
        RECT 113.165 55.715 113.335 55.885 ;
        RECT 113.625 55.715 113.795 55.885 ;
        RECT 114.085 55.715 114.255 55.885 ;
        RECT 114.545 55.715 114.715 55.885 ;
        RECT 115.005 55.715 115.175 55.885 ;
        RECT 115.465 55.715 115.635 55.885 ;
        RECT 115.925 55.715 116.095 55.885 ;
        RECT 116.385 55.715 116.555 55.885 ;
        RECT 116.845 55.715 117.015 55.885 ;
        RECT 117.305 55.715 117.475 55.885 ;
        RECT 117.765 55.715 117.935 55.885 ;
        RECT 118.225 55.715 118.395 55.885 ;
        RECT 118.685 55.715 118.855 55.885 ;
        RECT 119.145 55.715 119.315 55.885 ;
        RECT 119.605 55.715 119.775 55.885 ;
        RECT 120.065 55.715 120.235 55.885 ;
        RECT 120.525 55.715 120.695 55.885 ;
        RECT 120.985 55.715 121.155 55.885 ;
        RECT 121.445 55.715 121.615 55.885 ;
        RECT 121.905 55.715 122.075 55.885 ;
        RECT 122.365 55.715 122.535 55.885 ;
        RECT 122.825 55.715 122.995 55.885 ;
        RECT 123.285 55.715 123.455 55.885 ;
        RECT 123.745 55.715 123.915 55.885 ;
        RECT 124.205 55.715 124.375 55.885 ;
        RECT 124.665 55.715 124.835 55.885 ;
        RECT 125.125 55.715 125.295 55.885 ;
        RECT 125.585 55.715 125.755 55.885 ;
        RECT 126.045 55.715 126.215 55.885 ;
        RECT 126.505 55.715 126.675 55.885 ;
        RECT 126.965 55.715 127.135 55.885 ;
        RECT 127.425 55.715 127.595 55.885 ;
        RECT 127.885 55.715 128.055 55.885 ;
        RECT 128.345 55.715 128.515 55.885 ;
        RECT 128.805 55.715 128.975 55.885 ;
        RECT 129.265 55.715 129.435 55.885 ;
        RECT 129.725 55.715 129.895 55.885 ;
        RECT 130.185 55.715 130.355 55.885 ;
        RECT 130.645 55.715 130.815 55.885 ;
        RECT 131.105 55.715 131.275 55.885 ;
        RECT 131.565 55.715 131.735 55.885 ;
        RECT 132.025 55.715 132.195 55.885 ;
        RECT 132.485 55.715 132.655 55.885 ;
        RECT 132.945 55.715 133.115 55.885 ;
        RECT 133.405 55.715 133.575 55.885 ;
        RECT 133.865 55.715 134.035 55.885 ;
        RECT 134.325 55.715 134.495 55.885 ;
        RECT 134.785 55.715 134.955 55.885 ;
        RECT 135.245 55.715 135.415 55.885 ;
        RECT 135.705 55.715 135.875 55.885 ;
        RECT 136.165 55.715 136.335 55.885 ;
        RECT 136.625 55.715 136.795 55.885 ;
        RECT 137.085 55.715 137.255 55.885 ;
        RECT 137.545 55.715 137.715 55.885 ;
        RECT 138.005 55.715 138.175 55.885 ;
        RECT 138.465 55.715 138.635 55.885 ;
        RECT 138.925 55.715 139.095 55.885 ;
        RECT 139.385 55.715 139.555 55.885 ;
        RECT 139.845 55.715 140.015 55.885 ;
        RECT 140.305 55.715 140.475 55.885 ;
        RECT 140.765 55.715 140.935 55.885 ;
        RECT 141.225 55.715 141.395 55.885 ;
        RECT 141.685 55.715 141.855 55.885 ;
        RECT 142.145 55.715 142.315 55.885 ;
        RECT 142.605 55.715 142.775 55.885 ;
        RECT 143.065 55.715 143.235 55.885 ;
        RECT 143.525 55.715 143.695 55.885 ;
        RECT 143.985 55.715 144.155 55.885 ;
        RECT 55.665 50.275 55.835 50.445 ;
        RECT 56.125 50.275 56.295 50.445 ;
        RECT 56.585 50.275 56.755 50.445 ;
        RECT 57.045 50.275 57.215 50.445 ;
        RECT 57.505 50.275 57.675 50.445 ;
        RECT 57.965 50.275 58.135 50.445 ;
        RECT 58.425 50.275 58.595 50.445 ;
        RECT 58.885 50.275 59.055 50.445 ;
        RECT 59.345 50.275 59.515 50.445 ;
        RECT 59.805 50.275 59.975 50.445 ;
        RECT 60.265 50.275 60.435 50.445 ;
        RECT 60.725 50.275 60.895 50.445 ;
        RECT 61.185 50.275 61.355 50.445 ;
        RECT 61.645 50.275 61.815 50.445 ;
        RECT 62.105 50.275 62.275 50.445 ;
        RECT 62.565 50.275 62.735 50.445 ;
        RECT 63.025 50.275 63.195 50.445 ;
        RECT 63.485 50.275 63.655 50.445 ;
        RECT 63.945 50.275 64.115 50.445 ;
        RECT 64.405 50.275 64.575 50.445 ;
        RECT 64.865 50.275 65.035 50.445 ;
        RECT 65.325 50.275 65.495 50.445 ;
        RECT 65.785 50.275 65.955 50.445 ;
        RECT 66.245 50.275 66.415 50.445 ;
        RECT 66.705 50.275 66.875 50.445 ;
        RECT 67.165 50.275 67.335 50.445 ;
        RECT 67.625 50.275 67.795 50.445 ;
        RECT 68.085 50.275 68.255 50.445 ;
        RECT 68.545 50.275 68.715 50.445 ;
        RECT 69.005 50.275 69.175 50.445 ;
        RECT 69.465 50.275 69.635 50.445 ;
        RECT 69.925 50.275 70.095 50.445 ;
        RECT 70.385 50.275 70.555 50.445 ;
        RECT 70.845 50.275 71.015 50.445 ;
        RECT 71.305 50.275 71.475 50.445 ;
        RECT 71.765 50.275 71.935 50.445 ;
        RECT 72.225 50.275 72.395 50.445 ;
        RECT 72.685 50.275 72.855 50.445 ;
        RECT 73.145 50.275 73.315 50.445 ;
        RECT 73.605 50.275 73.775 50.445 ;
        RECT 74.065 50.275 74.235 50.445 ;
        RECT 74.525 50.275 74.695 50.445 ;
        RECT 74.985 50.275 75.155 50.445 ;
        RECT 75.445 50.275 75.615 50.445 ;
        RECT 75.905 50.275 76.075 50.445 ;
        RECT 76.365 50.275 76.535 50.445 ;
        RECT 76.825 50.275 76.995 50.445 ;
        RECT 77.285 50.275 77.455 50.445 ;
        RECT 77.745 50.275 77.915 50.445 ;
        RECT 78.205 50.275 78.375 50.445 ;
        RECT 78.665 50.275 78.835 50.445 ;
        RECT 79.125 50.275 79.295 50.445 ;
        RECT 79.585 50.275 79.755 50.445 ;
        RECT 80.045 50.275 80.215 50.445 ;
        RECT 80.505 50.275 80.675 50.445 ;
        RECT 80.965 50.275 81.135 50.445 ;
        RECT 81.425 50.275 81.595 50.445 ;
        RECT 81.885 50.275 82.055 50.445 ;
        RECT 82.345 50.275 82.515 50.445 ;
        RECT 82.805 50.275 82.975 50.445 ;
        RECT 83.265 50.275 83.435 50.445 ;
        RECT 83.725 50.275 83.895 50.445 ;
        RECT 84.185 50.275 84.355 50.445 ;
        RECT 84.645 50.275 84.815 50.445 ;
        RECT 85.105 50.275 85.275 50.445 ;
        RECT 85.565 50.275 85.735 50.445 ;
        RECT 86.025 50.275 86.195 50.445 ;
        RECT 86.485 50.275 86.655 50.445 ;
        RECT 86.945 50.275 87.115 50.445 ;
        RECT 87.405 50.275 87.575 50.445 ;
        RECT 87.865 50.275 88.035 50.445 ;
        RECT 88.325 50.275 88.495 50.445 ;
        RECT 88.785 50.275 88.955 50.445 ;
        RECT 89.245 50.275 89.415 50.445 ;
        RECT 89.705 50.275 89.875 50.445 ;
        RECT 90.165 50.275 90.335 50.445 ;
        RECT 90.625 50.275 90.795 50.445 ;
        RECT 91.085 50.275 91.255 50.445 ;
        RECT 91.545 50.275 91.715 50.445 ;
        RECT 92.005 50.275 92.175 50.445 ;
        RECT 92.465 50.275 92.635 50.445 ;
        RECT 92.925 50.275 93.095 50.445 ;
        RECT 93.385 50.275 93.555 50.445 ;
        RECT 93.845 50.275 94.015 50.445 ;
        RECT 94.305 50.275 94.475 50.445 ;
        RECT 94.765 50.275 94.935 50.445 ;
        RECT 95.225 50.275 95.395 50.445 ;
        RECT 95.685 50.275 95.855 50.445 ;
        RECT 96.145 50.275 96.315 50.445 ;
        RECT 96.605 50.275 96.775 50.445 ;
        RECT 97.065 50.275 97.235 50.445 ;
        RECT 97.525 50.275 97.695 50.445 ;
        RECT 97.985 50.275 98.155 50.445 ;
        RECT 98.445 50.275 98.615 50.445 ;
        RECT 98.905 50.275 99.075 50.445 ;
        RECT 99.365 50.275 99.535 50.445 ;
        RECT 99.825 50.275 99.995 50.445 ;
        RECT 100.285 50.275 100.455 50.445 ;
        RECT 100.745 50.275 100.915 50.445 ;
        RECT 101.205 50.275 101.375 50.445 ;
        RECT 101.665 50.275 101.835 50.445 ;
        RECT 102.125 50.275 102.295 50.445 ;
        RECT 102.585 50.275 102.755 50.445 ;
        RECT 103.045 50.275 103.215 50.445 ;
        RECT 103.505 50.275 103.675 50.445 ;
        RECT 103.965 50.275 104.135 50.445 ;
        RECT 104.425 50.275 104.595 50.445 ;
        RECT 104.885 50.275 105.055 50.445 ;
        RECT 105.345 50.275 105.515 50.445 ;
        RECT 105.805 50.275 105.975 50.445 ;
        RECT 106.265 50.275 106.435 50.445 ;
        RECT 106.725 50.275 106.895 50.445 ;
        RECT 107.185 50.275 107.355 50.445 ;
        RECT 107.645 50.275 107.815 50.445 ;
        RECT 108.105 50.275 108.275 50.445 ;
        RECT 108.565 50.275 108.735 50.445 ;
        RECT 109.025 50.275 109.195 50.445 ;
        RECT 109.485 50.275 109.655 50.445 ;
        RECT 109.945 50.275 110.115 50.445 ;
        RECT 110.405 50.275 110.575 50.445 ;
        RECT 110.865 50.275 111.035 50.445 ;
        RECT 111.325 50.275 111.495 50.445 ;
        RECT 111.785 50.275 111.955 50.445 ;
        RECT 112.245 50.275 112.415 50.445 ;
        RECT 112.705 50.275 112.875 50.445 ;
        RECT 113.165 50.275 113.335 50.445 ;
        RECT 113.625 50.275 113.795 50.445 ;
        RECT 114.085 50.275 114.255 50.445 ;
        RECT 114.545 50.275 114.715 50.445 ;
        RECT 115.005 50.275 115.175 50.445 ;
        RECT 115.465 50.275 115.635 50.445 ;
        RECT 115.925 50.275 116.095 50.445 ;
        RECT 116.385 50.275 116.555 50.445 ;
        RECT 116.845 50.275 117.015 50.445 ;
        RECT 117.305 50.275 117.475 50.445 ;
        RECT 117.765 50.275 117.935 50.445 ;
        RECT 118.225 50.275 118.395 50.445 ;
        RECT 118.685 50.275 118.855 50.445 ;
        RECT 119.145 50.275 119.315 50.445 ;
        RECT 119.605 50.275 119.775 50.445 ;
        RECT 120.065 50.275 120.235 50.445 ;
        RECT 120.525 50.275 120.695 50.445 ;
        RECT 120.985 50.275 121.155 50.445 ;
        RECT 121.445 50.275 121.615 50.445 ;
        RECT 121.905 50.275 122.075 50.445 ;
        RECT 122.365 50.275 122.535 50.445 ;
        RECT 122.825 50.275 122.995 50.445 ;
        RECT 123.285 50.275 123.455 50.445 ;
        RECT 123.745 50.275 123.915 50.445 ;
        RECT 124.205 50.275 124.375 50.445 ;
        RECT 124.665 50.275 124.835 50.445 ;
        RECT 125.125 50.275 125.295 50.445 ;
        RECT 125.585 50.275 125.755 50.445 ;
        RECT 126.045 50.275 126.215 50.445 ;
        RECT 126.505 50.275 126.675 50.445 ;
        RECT 126.965 50.275 127.135 50.445 ;
        RECT 127.425 50.275 127.595 50.445 ;
        RECT 127.885 50.275 128.055 50.445 ;
        RECT 128.345 50.275 128.515 50.445 ;
        RECT 128.805 50.275 128.975 50.445 ;
        RECT 129.265 50.275 129.435 50.445 ;
        RECT 129.725 50.275 129.895 50.445 ;
        RECT 130.185 50.275 130.355 50.445 ;
        RECT 130.645 50.275 130.815 50.445 ;
        RECT 131.105 50.275 131.275 50.445 ;
        RECT 131.565 50.275 131.735 50.445 ;
        RECT 132.025 50.275 132.195 50.445 ;
        RECT 132.485 50.275 132.655 50.445 ;
        RECT 132.945 50.275 133.115 50.445 ;
        RECT 133.405 50.275 133.575 50.445 ;
        RECT 133.865 50.275 134.035 50.445 ;
        RECT 134.325 50.275 134.495 50.445 ;
        RECT 134.785 50.275 134.955 50.445 ;
        RECT 135.245 50.275 135.415 50.445 ;
        RECT 135.705 50.275 135.875 50.445 ;
        RECT 136.165 50.275 136.335 50.445 ;
        RECT 136.625 50.275 136.795 50.445 ;
        RECT 137.085 50.275 137.255 50.445 ;
        RECT 137.545 50.275 137.715 50.445 ;
        RECT 138.005 50.275 138.175 50.445 ;
        RECT 138.465 50.275 138.635 50.445 ;
        RECT 138.925 50.275 139.095 50.445 ;
        RECT 139.385 50.275 139.555 50.445 ;
        RECT 139.845 50.275 140.015 50.445 ;
        RECT 140.305 50.275 140.475 50.445 ;
        RECT 140.765 50.275 140.935 50.445 ;
        RECT 141.225 50.275 141.395 50.445 ;
        RECT 141.685 50.275 141.855 50.445 ;
        RECT 142.145 50.275 142.315 50.445 ;
        RECT 142.605 50.275 142.775 50.445 ;
        RECT 143.065 50.275 143.235 50.445 ;
        RECT 143.525 50.275 143.695 50.445 ;
        RECT 143.985 50.275 144.155 50.445 ;
        RECT 55.665 44.835 55.835 45.005 ;
        RECT 56.125 44.835 56.295 45.005 ;
        RECT 56.585 44.835 56.755 45.005 ;
        RECT 57.045 44.835 57.215 45.005 ;
        RECT 57.505 44.835 57.675 45.005 ;
        RECT 57.965 44.835 58.135 45.005 ;
        RECT 58.425 44.835 58.595 45.005 ;
        RECT 58.885 44.835 59.055 45.005 ;
        RECT 59.345 44.835 59.515 45.005 ;
        RECT 59.805 44.835 59.975 45.005 ;
        RECT 60.265 44.835 60.435 45.005 ;
        RECT 60.725 44.835 60.895 45.005 ;
        RECT 61.185 44.835 61.355 45.005 ;
        RECT 61.645 44.835 61.815 45.005 ;
        RECT 62.105 44.835 62.275 45.005 ;
        RECT 62.565 44.835 62.735 45.005 ;
        RECT 63.025 44.835 63.195 45.005 ;
        RECT 63.485 44.835 63.655 45.005 ;
        RECT 63.945 44.835 64.115 45.005 ;
        RECT 64.405 44.835 64.575 45.005 ;
        RECT 64.865 44.835 65.035 45.005 ;
        RECT 65.325 44.835 65.495 45.005 ;
        RECT 65.785 44.835 65.955 45.005 ;
        RECT 66.245 44.835 66.415 45.005 ;
        RECT 66.705 44.835 66.875 45.005 ;
        RECT 67.165 44.835 67.335 45.005 ;
        RECT 67.625 44.835 67.795 45.005 ;
        RECT 68.085 44.835 68.255 45.005 ;
        RECT 68.545 44.835 68.715 45.005 ;
        RECT 69.005 44.835 69.175 45.005 ;
        RECT 69.465 44.835 69.635 45.005 ;
        RECT 69.925 44.835 70.095 45.005 ;
        RECT 70.385 44.835 70.555 45.005 ;
        RECT 70.845 44.835 71.015 45.005 ;
        RECT 71.305 44.835 71.475 45.005 ;
        RECT 71.765 44.835 71.935 45.005 ;
        RECT 72.225 44.835 72.395 45.005 ;
        RECT 72.685 44.835 72.855 45.005 ;
        RECT 73.145 44.835 73.315 45.005 ;
        RECT 73.605 44.835 73.775 45.005 ;
        RECT 74.065 44.835 74.235 45.005 ;
        RECT 74.525 44.835 74.695 45.005 ;
        RECT 74.985 44.835 75.155 45.005 ;
        RECT 75.445 44.835 75.615 45.005 ;
        RECT 75.905 44.835 76.075 45.005 ;
        RECT 76.365 44.835 76.535 45.005 ;
        RECT 76.825 44.835 76.995 45.005 ;
        RECT 77.285 44.835 77.455 45.005 ;
        RECT 77.745 44.835 77.915 45.005 ;
        RECT 78.205 44.835 78.375 45.005 ;
        RECT 78.665 44.835 78.835 45.005 ;
        RECT 79.125 44.835 79.295 45.005 ;
        RECT 79.585 44.835 79.755 45.005 ;
        RECT 80.045 44.835 80.215 45.005 ;
        RECT 80.505 44.835 80.675 45.005 ;
        RECT 80.965 44.835 81.135 45.005 ;
        RECT 81.425 44.835 81.595 45.005 ;
        RECT 81.885 44.835 82.055 45.005 ;
        RECT 82.345 44.835 82.515 45.005 ;
        RECT 82.805 44.835 82.975 45.005 ;
        RECT 83.265 44.835 83.435 45.005 ;
        RECT 83.725 44.835 83.895 45.005 ;
        RECT 84.185 44.835 84.355 45.005 ;
        RECT 84.645 44.835 84.815 45.005 ;
        RECT 85.105 44.835 85.275 45.005 ;
        RECT 85.565 44.835 85.735 45.005 ;
        RECT 86.025 44.835 86.195 45.005 ;
        RECT 86.485 44.835 86.655 45.005 ;
        RECT 86.945 44.835 87.115 45.005 ;
        RECT 87.405 44.835 87.575 45.005 ;
        RECT 87.865 44.835 88.035 45.005 ;
        RECT 88.325 44.835 88.495 45.005 ;
        RECT 88.785 44.835 88.955 45.005 ;
        RECT 89.245 44.835 89.415 45.005 ;
        RECT 89.705 44.835 89.875 45.005 ;
        RECT 90.165 44.835 90.335 45.005 ;
        RECT 90.625 44.835 90.795 45.005 ;
        RECT 91.085 44.835 91.255 45.005 ;
        RECT 91.545 44.835 91.715 45.005 ;
        RECT 92.005 44.835 92.175 45.005 ;
        RECT 92.465 44.835 92.635 45.005 ;
        RECT 92.925 44.835 93.095 45.005 ;
        RECT 93.385 44.835 93.555 45.005 ;
        RECT 93.845 44.835 94.015 45.005 ;
        RECT 94.305 44.835 94.475 45.005 ;
        RECT 94.765 44.835 94.935 45.005 ;
        RECT 95.225 44.835 95.395 45.005 ;
        RECT 95.685 44.835 95.855 45.005 ;
        RECT 96.145 44.835 96.315 45.005 ;
        RECT 96.605 44.835 96.775 45.005 ;
        RECT 97.065 44.835 97.235 45.005 ;
        RECT 97.525 44.835 97.695 45.005 ;
        RECT 97.985 44.835 98.155 45.005 ;
        RECT 98.445 44.835 98.615 45.005 ;
        RECT 98.905 44.835 99.075 45.005 ;
        RECT 99.365 44.835 99.535 45.005 ;
        RECT 99.825 44.835 99.995 45.005 ;
        RECT 100.285 44.835 100.455 45.005 ;
        RECT 100.745 44.835 100.915 45.005 ;
        RECT 101.205 44.835 101.375 45.005 ;
        RECT 101.665 44.835 101.835 45.005 ;
        RECT 102.125 44.835 102.295 45.005 ;
        RECT 102.585 44.835 102.755 45.005 ;
        RECT 103.045 44.835 103.215 45.005 ;
        RECT 103.505 44.835 103.675 45.005 ;
        RECT 103.965 44.835 104.135 45.005 ;
        RECT 104.425 44.835 104.595 45.005 ;
        RECT 104.885 44.835 105.055 45.005 ;
        RECT 105.345 44.835 105.515 45.005 ;
        RECT 105.805 44.835 105.975 45.005 ;
        RECT 106.265 44.835 106.435 45.005 ;
        RECT 106.725 44.835 106.895 45.005 ;
        RECT 107.185 44.835 107.355 45.005 ;
        RECT 107.645 44.835 107.815 45.005 ;
        RECT 108.105 44.835 108.275 45.005 ;
        RECT 108.565 44.835 108.735 45.005 ;
        RECT 109.025 44.835 109.195 45.005 ;
        RECT 109.485 44.835 109.655 45.005 ;
        RECT 109.945 44.835 110.115 45.005 ;
        RECT 110.405 44.835 110.575 45.005 ;
        RECT 110.865 44.835 111.035 45.005 ;
        RECT 111.325 44.835 111.495 45.005 ;
        RECT 111.785 44.835 111.955 45.005 ;
        RECT 112.245 44.835 112.415 45.005 ;
        RECT 112.705 44.835 112.875 45.005 ;
        RECT 113.165 44.835 113.335 45.005 ;
        RECT 113.625 44.835 113.795 45.005 ;
        RECT 114.085 44.835 114.255 45.005 ;
        RECT 114.545 44.835 114.715 45.005 ;
        RECT 115.005 44.835 115.175 45.005 ;
        RECT 115.465 44.835 115.635 45.005 ;
        RECT 115.925 44.835 116.095 45.005 ;
        RECT 116.385 44.835 116.555 45.005 ;
        RECT 116.845 44.835 117.015 45.005 ;
        RECT 117.305 44.835 117.475 45.005 ;
        RECT 117.765 44.835 117.935 45.005 ;
        RECT 118.225 44.835 118.395 45.005 ;
        RECT 118.685 44.835 118.855 45.005 ;
        RECT 119.145 44.835 119.315 45.005 ;
        RECT 119.605 44.835 119.775 45.005 ;
        RECT 120.065 44.835 120.235 45.005 ;
        RECT 120.525 44.835 120.695 45.005 ;
        RECT 120.985 44.835 121.155 45.005 ;
        RECT 121.445 44.835 121.615 45.005 ;
        RECT 121.905 44.835 122.075 45.005 ;
        RECT 122.365 44.835 122.535 45.005 ;
        RECT 122.825 44.835 122.995 45.005 ;
        RECT 123.285 44.835 123.455 45.005 ;
        RECT 123.745 44.835 123.915 45.005 ;
        RECT 124.205 44.835 124.375 45.005 ;
        RECT 124.665 44.835 124.835 45.005 ;
        RECT 125.125 44.835 125.295 45.005 ;
        RECT 125.585 44.835 125.755 45.005 ;
        RECT 126.045 44.835 126.215 45.005 ;
        RECT 126.505 44.835 126.675 45.005 ;
        RECT 126.965 44.835 127.135 45.005 ;
        RECT 127.425 44.835 127.595 45.005 ;
        RECT 127.885 44.835 128.055 45.005 ;
        RECT 128.345 44.835 128.515 45.005 ;
        RECT 128.805 44.835 128.975 45.005 ;
        RECT 129.265 44.835 129.435 45.005 ;
        RECT 129.725 44.835 129.895 45.005 ;
        RECT 130.185 44.835 130.355 45.005 ;
        RECT 130.645 44.835 130.815 45.005 ;
        RECT 131.105 44.835 131.275 45.005 ;
        RECT 131.565 44.835 131.735 45.005 ;
        RECT 132.025 44.835 132.195 45.005 ;
        RECT 132.485 44.835 132.655 45.005 ;
        RECT 132.945 44.835 133.115 45.005 ;
        RECT 133.405 44.835 133.575 45.005 ;
        RECT 133.865 44.835 134.035 45.005 ;
        RECT 134.325 44.835 134.495 45.005 ;
        RECT 134.785 44.835 134.955 45.005 ;
        RECT 135.245 44.835 135.415 45.005 ;
        RECT 135.705 44.835 135.875 45.005 ;
        RECT 136.165 44.835 136.335 45.005 ;
        RECT 136.625 44.835 136.795 45.005 ;
        RECT 137.085 44.835 137.255 45.005 ;
        RECT 137.545 44.835 137.715 45.005 ;
        RECT 138.005 44.835 138.175 45.005 ;
        RECT 138.465 44.835 138.635 45.005 ;
        RECT 138.925 44.835 139.095 45.005 ;
        RECT 139.385 44.835 139.555 45.005 ;
        RECT 139.845 44.835 140.015 45.005 ;
        RECT 140.305 44.835 140.475 45.005 ;
        RECT 140.765 44.835 140.935 45.005 ;
        RECT 141.225 44.835 141.395 45.005 ;
        RECT 141.685 44.835 141.855 45.005 ;
        RECT 142.145 44.835 142.315 45.005 ;
        RECT 142.605 44.835 142.775 45.005 ;
        RECT 143.065 44.835 143.235 45.005 ;
        RECT 143.525 44.835 143.695 45.005 ;
        RECT 143.985 44.835 144.155 45.005 ;
        RECT 55.665 39.395 55.835 39.565 ;
        RECT 56.125 39.395 56.295 39.565 ;
        RECT 56.585 39.395 56.755 39.565 ;
        RECT 57.045 39.395 57.215 39.565 ;
        RECT 57.505 39.395 57.675 39.565 ;
        RECT 57.965 39.395 58.135 39.565 ;
        RECT 58.425 39.395 58.595 39.565 ;
        RECT 58.885 39.395 59.055 39.565 ;
        RECT 59.345 39.395 59.515 39.565 ;
        RECT 59.805 39.395 59.975 39.565 ;
        RECT 60.265 39.395 60.435 39.565 ;
        RECT 60.725 39.395 60.895 39.565 ;
        RECT 61.185 39.395 61.355 39.565 ;
        RECT 61.645 39.395 61.815 39.565 ;
        RECT 62.105 39.395 62.275 39.565 ;
        RECT 62.565 39.395 62.735 39.565 ;
        RECT 63.025 39.395 63.195 39.565 ;
        RECT 63.485 39.395 63.655 39.565 ;
        RECT 63.945 39.395 64.115 39.565 ;
        RECT 64.405 39.395 64.575 39.565 ;
        RECT 64.865 39.395 65.035 39.565 ;
        RECT 65.325 39.395 65.495 39.565 ;
        RECT 65.785 39.395 65.955 39.565 ;
        RECT 66.245 39.395 66.415 39.565 ;
        RECT 66.705 39.395 66.875 39.565 ;
        RECT 67.165 39.395 67.335 39.565 ;
        RECT 67.625 39.395 67.795 39.565 ;
        RECT 68.085 39.395 68.255 39.565 ;
        RECT 68.545 39.395 68.715 39.565 ;
        RECT 69.005 39.395 69.175 39.565 ;
        RECT 69.465 39.395 69.635 39.565 ;
        RECT 69.925 39.395 70.095 39.565 ;
        RECT 70.385 39.395 70.555 39.565 ;
        RECT 70.845 39.395 71.015 39.565 ;
        RECT 71.305 39.395 71.475 39.565 ;
        RECT 71.765 39.395 71.935 39.565 ;
        RECT 72.225 39.395 72.395 39.565 ;
        RECT 72.685 39.395 72.855 39.565 ;
        RECT 73.145 39.395 73.315 39.565 ;
        RECT 73.605 39.395 73.775 39.565 ;
        RECT 74.065 39.395 74.235 39.565 ;
        RECT 74.525 39.395 74.695 39.565 ;
        RECT 74.985 39.395 75.155 39.565 ;
        RECT 75.445 39.395 75.615 39.565 ;
        RECT 75.905 39.395 76.075 39.565 ;
        RECT 76.365 39.395 76.535 39.565 ;
        RECT 76.825 39.395 76.995 39.565 ;
        RECT 77.285 39.395 77.455 39.565 ;
        RECT 77.745 39.395 77.915 39.565 ;
        RECT 78.205 39.395 78.375 39.565 ;
        RECT 78.665 39.395 78.835 39.565 ;
        RECT 79.125 39.395 79.295 39.565 ;
        RECT 79.585 39.395 79.755 39.565 ;
        RECT 80.045 39.395 80.215 39.565 ;
        RECT 80.505 39.395 80.675 39.565 ;
        RECT 80.965 39.395 81.135 39.565 ;
        RECT 81.425 39.395 81.595 39.565 ;
        RECT 81.885 39.395 82.055 39.565 ;
        RECT 82.345 39.395 82.515 39.565 ;
        RECT 82.805 39.395 82.975 39.565 ;
        RECT 83.265 39.395 83.435 39.565 ;
        RECT 83.725 39.395 83.895 39.565 ;
        RECT 84.185 39.395 84.355 39.565 ;
        RECT 84.645 39.395 84.815 39.565 ;
        RECT 85.105 39.395 85.275 39.565 ;
        RECT 85.565 39.395 85.735 39.565 ;
        RECT 86.025 39.395 86.195 39.565 ;
        RECT 86.485 39.395 86.655 39.565 ;
        RECT 86.945 39.395 87.115 39.565 ;
        RECT 87.405 39.395 87.575 39.565 ;
        RECT 87.865 39.395 88.035 39.565 ;
        RECT 88.325 39.395 88.495 39.565 ;
        RECT 88.785 39.395 88.955 39.565 ;
        RECT 89.245 39.395 89.415 39.565 ;
        RECT 89.705 39.395 89.875 39.565 ;
        RECT 90.165 39.395 90.335 39.565 ;
        RECT 90.625 39.395 90.795 39.565 ;
        RECT 91.085 39.395 91.255 39.565 ;
        RECT 91.545 39.395 91.715 39.565 ;
        RECT 92.005 39.395 92.175 39.565 ;
        RECT 92.465 39.395 92.635 39.565 ;
        RECT 92.925 39.395 93.095 39.565 ;
        RECT 93.385 39.395 93.555 39.565 ;
        RECT 93.845 39.395 94.015 39.565 ;
        RECT 94.305 39.395 94.475 39.565 ;
        RECT 94.765 39.395 94.935 39.565 ;
        RECT 95.225 39.395 95.395 39.565 ;
        RECT 95.685 39.395 95.855 39.565 ;
        RECT 96.145 39.395 96.315 39.565 ;
        RECT 96.605 39.395 96.775 39.565 ;
        RECT 97.065 39.395 97.235 39.565 ;
        RECT 97.525 39.395 97.695 39.565 ;
        RECT 97.985 39.395 98.155 39.565 ;
        RECT 98.445 39.395 98.615 39.565 ;
        RECT 98.905 39.395 99.075 39.565 ;
        RECT 99.365 39.395 99.535 39.565 ;
        RECT 99.825 39.395 99.995 39.565 ;
        RECT 100.285 39.395 100.455 39.565 ;
        RECT 100.745 39.395 100.915 39.565 ;
        RECT 101.205 39.395 101.375 39.565 ;
        RECT 101.665 39.395 101.835 39.565 ;
        RECT 102.125 39.395 102.295 39.565 ;
        RECT 102.585 39.395 102.755 39.565 ;
        RECT 103.045 39.395 103.215 39.565 ;
        RECT 103.505 39.395 103.675 39.565 ;
        RECT 103.965 39.395 104.135 39.565 ;
        RECT 104.425 39.395 104.595 39.565 ;
        RECT 104.885 39.395 105.055 39.565 ;
        RECT 105.345 39.395 105.515 39.565 ;
        RECT 105.805 39.395 105.975 39.565 ;
        RECT 106.265 39.395 106.435 39.565 ;
        RECT 106.725 39.395 106.895 39.565 ;
        RECT 107.185 39.395 107.355 39.565 ;
        RECT 107.645 39.395 107.815 39.565 ;
        RECT 108.105 39.395 108.275 39.565 ;
        RECT 108.565 39.395 108.735 39.565 ;
        RECT 109.025 39.395 109.195 39.565 ;
        RECT 109.485 39.395 109.655 39.565 ;
        RECT 109.945 39.395 110.115 39.565 ;
        RECT 110.405 39.395 110.575 39.565 ;
        RECT 110.865 39.395 111.035 39.565 ;
        RECT 111.325 39.395 111.495 39.565 ;
        RECT 111.785 39.395 111.955 39.565 ;
        RECT 112.245 39.395 112.415 39.565 ;
        RECT 112.705 39.395 112.875 39.565 ;
        RECT 113.165 39.395 113.335 39.565 ;
        RECT 113.625 39.395 113.795 39.565 ;
        RECT 114.085 39.395 114.255 39.565 ;
        RECT 114.545 39.395 114.715 39.565 ;
        RECT 115.005 39.395 115.175 39.565 ;
        RECT 115.465 39.395 115.635 39.565 ;
        RECT 115.925 39.395 116.095 39.565 ;
        RECT 116.385 39.395 116.555 39.565 ;
        RECT 116.845 39.395 117.015 39.565 ;
        RECT 117.305 39.395 117.475 39.565 ;
        RECT 117.765 39.395 117.935 39.565 ;
        RECT 118.225 39.395 118.395 39.565 ;
        RECT 118.685 39.395 118.855 39.565 ;
        RECT 119.145 39.395 119.315 39.565 ;
        RECT 119.605 39.395 119.775 39.565 ;
        RECT 120.065 39.395 120.235 39.565 ;
        RECT 120.525 39.395 120.695 39.565 ;
        RECT 120.985 39.395 121.155 39.565 ;
        RECT 121.445 39.395 121.615 39.565 ;
        RECT 121.905 39.395 122.075 39.565 ;
        RECT 122.365 39.395 122.535 39.565 ;
        RECT 122.825 39.395 122.995 39.565 ;
        RECT 123.285 39.395 123.455 39.565 ;
        RECT 123.745 39.395 123.915 39.565 ;
        RECT 124.205 39.395 124.375 39.565 ;
        RECT 124.665 39.395 124.835 39.565 ;
        RECT 125.125 39.395 125.295 39.565 ;
        RECT 125.585 39.395 125.755 39.565 ;
        RECT 126.045 39.395 126.215 39.565 ;
        RECT 126.505 39.395 126.675 39.565 ;
        RECT 126.965 39.395 127.135 39.565 ;
        RECT 127.425 39.395 127.595 39.565 ;
        RECT 127.885 39.395 128.055 39.565 ;
        RECT 128.345 39.395 128.515 39.565 ;
        RECT 128.805 39.395 128.975 39.565 ;
        RECT 129.265 39.395 129.435 39.565 ;
        RECT 129.725 39.395 129.895 39.565 ;
        RECT 130.185 39.395 130.355 39.565 ;
        RECT 130.645 39.395 130.815 39.565 ;
        RECT 131.105 39.395 131.275 39.565 ;
        RECT 131.565 39.395 131.735 39.565 ;
        RECT 132.025 39.395 132.195 39.565 ;
        RECT 132.485 39.395 132.655 39.565 ;
        RECT 132.945 39.395 133.115 39.565 ;
        RECT 133.405 39.395 133.575 39.565 ;
        RECT 133.865 39.395 134.035 39.565 ;
        RECT 134.325 39.395 134.495 39.565 ;
        RECT 134.785 39.395 134.955 39.565 ;
        RECT 135.245 39.395 135.415 39.565 ;
        RECT 135.705 39.395 135.875 39.565 ;
        RECT 136.165 39.395 136.335 39.565 ;
        RECT 136.625 39.395 136.795 39.565 ;
        RECT 137.085 39.395 137.255 39.565 ;
        RECT 137.545 39.395 137.715 39.565 ;
        RECT 138.005 39.395 138.175 39.565 ;
        RECT 138.465 39.395 138.635 39.565 ;
        RECT 138.925 39.395 139.095 39.565 ;
        RECT 139.385 39.395 139.555 39.565 ;
        RECT 139.845 39.395 140.015 39.565 ;
        RECT 140.305 39.395 140.475 39.565 ;
        RECT 140.765 39.395 140.935 39.565 ;
        RECT 141.225 39.395 141.395 39.565 ;
        RECT 141.685 39.395 141.855 39.565 ;
        RECT 142.145 39.395 142.315 39.565 ;
        RECT 142.605 39.395 142.775 39.565 ;
        RECT 143.065 39.395 143.235 39.565 ;
        RECT 143.525 39.395 143.695 39.565 ;
        RECT 143.985 39.395 144.155 39.565 ;
        RECT 55.665 33.955 55.835 34.125 ;
        RECT 56.125 33.955 56.295 34.125 ;
        RECT 56.585 33.955 56.755 34.125 ;
        RECT 57.045 33.955 57.215 34.125 ;
        RECT 57.505 33.955 57.675 34.125 ;
        RECT 57.965 33.955 58.135 34.125 ;
        RECT 58.425 33.955 58.595 34.125 ;
        RECT 58.885 33.955 59.055 34.125 ;
        RECT 59.345 33.955 59.515 34.125 ;
        RECT 59.805 33.955 59.975 34.125 ;
        RECT 60.265 33.955 60.435 34.125 ;
        RECT 60.725 33.955 60.895 34.125 ;
        RECT 61.185 33.955 61.355 34.125 ;
        RECT 61.645 33.955 61.815 34.125 ;
        RECT 62.105 33.955 62.275 34.125 ;
        RECT 62.565 33.955 62.735 34.125 ;
        RECT 63.025 33.955 63.195 34.125 ;
        RECT 63.485 33.955 63.655 34.125 ;
        RECT 63.945 33.955 64.115 34.125 ;
        RECT 64.405 33.955 64.575 34.125 ;
        RECT 64.865 33.955 65.035 34.125 ;
        RECT 65.325 33.955 65.495 34.125 ;
        RECT 65.785 33.955 65.955 34.125 ;
        RECT 66.245 33.955 66.415 34.125 ;
        RECT 66.705 33.955 66.875 34.125 ;
        RECT 67.165 33.955 67.335 34.125 ;
        RECT 67.625 33.955 67.795 34.125 ;
        RECT 68.085 33.955 68.255 34.125 ;
        RECT 68.545 33.955 68.715 34.125 ;
        RECT 69.005 33.955 69.175 34.125 ;
        RECT 69.465 33.955 69.635 34.125 ;
        RECT 69.925 33.955 70.095 34.125 ;
        RECT 70.385 33.955 70.555 34.125 ;
        RECT 70.845 33.955 71.015 34.125 ;
        RECT 71.305 33.955 71.475 34.125 ;
        RECT 71.765 33.955 71.935 34.125 ;
        RECT 72.225 33.955 72.395 34.125 ;
        RECT 72.685 33.955 72.855 34.125 ;
        RECT 73.145 33.955 73.315 34.125 ;
        RECT 73.605 33.955 73.775 34.125 ;
        RECT 74.065 33.955 74.235 34.125 ;
        RECT 74.525 33.955 74.695 34.125 ;
        RECT 74.985 33.955 75.155 34.125 ;
        RECT 75.445 33.955 75.615 34.125 ;
        RECT 75.905 33.955 76.075 34.125 ;
        RECT 76.365 33.955 76.535 34.125 ;
        RECT 76.825 33.955 76.995 34.125 ;
        RECT 77.285 33.955 77.455 34.125 ;
        RECT 77.745 33.955 77.915 34.125 ;
        RECT 78.205 33.955 78.375 34.125 ;
        RECT 78.665 33.955 78.835 34.125 ;
        RECT 79.125 33.955 79.295 34.125 ;
        RECT 79.585 33.955 79.755 34.125 ;
        RECT 80.045 33.955 80.215 34.125 ;
        RECT 80.505 33.955 80.675 34.125 ;
        RECT 80.965 33.955 81.135 34.125 ;
        RECT 81.425 33.955 81.595 34.125 ;
        RECT 81.885 33.955 82.055 34.125 ;
        RECT 82.345 33.955 82.515 34.125 ;
        RECT 82.805 33.955 82.975 34.125 ;
        RECT 83.265 33.955 83.435 34.125 ;
        RECT 83.725 33.955 83.895 34.125 ;
        RECT 84.185 33.955 84.355 34.125 ;
        RECT 84.645 33.955 84.815 34.125 ;
        RECT 85.105 33.955 85.275 34.125 ;
        RECT 85.565 33.955 85.735 34.125 ;
        RECT 86.025 33.955 86.195 34.125 ;
        RECT 86.485 33.955 86.655 34.125 ;
        RECT 86.945 33.955 87.115 34.125 ;
        RECT 87.405 33.955 87.575 34.125 ;
        RECT 87.865 33.955 88.035 34.125 ;
        RECT 88.325 33.955 88.495 34.125 ;
        RECT 88.785 33.955 88.955 34.125 ;
        RECT 89.245 33.955 89.415 34.125 ;
        RECT 89.705 33.955 89.875 34.125 ;
        RECT 90.165 33.955 90.335 34.125 ;
        RECT 90.625 33.955 90.795 34.125 ;
        RECT 91.085 33.955 91.255 34.125 ;
        RECT 91.545 33.955 91.715 34.125 ;
        RECT 92.005 33.955 92.175 34.125 ;
        RECT 92.465 33.955 92.635 34.125 ;
        RECT 92.925 33.955 93.095 34.125 ;
        RECT 93.385 33.955 93.555 34.125 ;
        RECT 93.845 33.955 94.015 34.125 ;
        RECT 94.305 33.955 94.475 34.125 ;
        RECT 94.765 33.955 94.935 34.125 ;
        RECT 95.225 33.955 95.395 34.125 ;
        RECT 95.685 33.955 95.855 34.125 ;
        RECT 96.145 33.955 96.315 34.125 ;
        RECT 96.605 33.955 96.775 34.125 ;
        RECT 97.065 33.955 97.235 34.125 ;
        RECT 97.525 33.955 97.695 34.125 ;
        RECT 97.985 33.955 98.155 34.125 ;
        RECT 98.445 33.955 98.615 34.125 ;
        RECT 98.905 33.955 99.075 34.125 ;
        RECT 99.365 33.955 99.535 34.125 ;
        RECT 99.825 33.955 99.995 34.125 ;
        RECT 100.285 33.955 100.455 34.125 ;
        RECT 100.745 33.955 100.915 34.125 ;
        RECT 101.205 33.955 101.375 34.125 ;
        RECT 101.665 33.955 101.835 34.125 ;
        RECT 102.125 33.955 102.295 34.125 ;
        RECT 102.585 33.955 102.755 34.125 ;
        RECT 103.045 33.955 103.215 34.125 ;
        RECT 103.505 33.955 103.675 34.125 ;
        RECT 103.965 33.955 104.135 34.125 ;
        RECT 104.425 33.955 104.595 34.125 ;
        RECT 104.885 33.955 105.055 34.125 ;
        RECT 105.345 33.955 105.515 34.125 ;
        RECT 105.805 33.955 105.975 34.125 ;
        RECT 106.265 33.955 106.435 34.125 ;
        RECT 106.725 33.955 106.895 34.125 ;
        RECT 107.185 33.955 107.355 34.125 ;
        RECT 107.645 33.955 107.815 34.125 ;
        RECT 108.105 33.955 108.275 34.125 ;
        RECT 108.565 33.955 108.735 34.125 ;
        RECT 109.025 33.955 109.195 34.125 ;
        RECT 109.485 33.955 109.655 34.125 ;
        RECT 109.945 33.955 110.115 34.125 ;
        RECT 110.405 33.955 110.575 34.125 ;
        RECT 110.865 33.955 111.035 34.125 ;
        RECT 111.325 33.955 111.495 34.125 ;
        RECT 111.785 33.955 111.955 34.125 ;
        RECT 112.245 33.955 112.415 34.125 ;
        RECT 112.705 33.955 112.875 34.125 ;
        RECT 113.165 33.955 113.335 34.125 ;
        RECT 113.625 33.955 113.795 34.125 ;
        RECT 114.085 33.955 114.255 34.125 ;
        RECT 114.545 33.955 114.715 34.125 ;
        RECT 115.005 33.955 115.175 34.125 ;
        RECT 115.465 33.955 115.635 34.125 ;
        RECT 115.925 33.955 116.095 34.125 ;
        RECT 116.385 33.955 116.555 34.125 ;
        RECT 116.845 33.955 117.015 34.125 ;
        RECT 117.305 33.955 117.475 34.125 ;
        RECT 117.765 33.955 117.935 34.125 ;
        RECT 118.225 33.955 118.395 34.125 ;
        RECT 118.685 33.955 118.855 34.125 ;
        RECT 119.145 33.955 119.315 34.125 ;
        RECT 119.605 33.955 119.775 34.125 ;
        RECT 120.065 33.955 120.235 34.125 ;
        RECT 120.525 33.955 120.695 34.125 ;
        RECT 120.985 33.955 121.155 34.125 ;
        RECT 121.445 33.955 121.615 34.125 ;
        RECT 121.905 33.955 122.075 34.125 ;
        RECT 122.365 33.955 122.535 34.125 ;
        RECT 122.825 33.955 122.995 34.125 ;
        RECT 123.285 33.955 123.455 34.125 ;
        RECT 123.745 33.955 123.915 34.125 ;
        RECT 124.205 33.955 124.375 34.125 ;
        RECT 124.665 33.955 124.835 34.125 ;
        RECT 125.125 33.955 125.295 34.125 ;
        RECT 125.585 33.955 125.755 34.125 ;
        RECT 126.045 33.955 126.215 34.125 ;
        RECT 126.505 33.955 126.675 34.125 ;
        RECT 126.965 33.955 127.135 34.125 ;
        RECT 127.425 33.955 127.595 34.125 ;
        RECT 127.885 33.955 128.055 34.125 ;
        RECT 128.345 33.955 128.515 34.125 ;
        RECT 128.805 33.955 128.975 34.125 ;
        RECT 129.265 33.955 129.435 34.125 ;
        RECT 129.725 33.955 129.895 34.125 ;
        RECT 130.185 33.955 130.355 34.125 ;
        RECT 130.645 33.955 130.815 34.125 ;
        RECT 131.105 33.955 131.275 34.125 ;
        RECT 131.565 33.955 131.735 34.125 ;
        RECT 132.025 33.955 132.195 34.125 ;
        RECT 132.485 33.955 132.655 34.125 ;
        RECT 132.945 33.955 133.115 34.125 ;
        RECT 133.405 33.955 133.575 34.125 ;
        RECT 133.865 33.955 134.035 34.125 ;
        RECT 134.325 33.955 134.495 34.125 ;
        RECT 134.785 33.955 134.955 34.125 ;
        RECT 135.245 33.955 135.415 34.125 ;
        RECT 135.705 33.955 135.875 34.125 ;
        RECT 136.165 33.955 136.335 34.125 ;
        RECT 136.625 33.955 136.795 34.125 ;
        RECT 137.085 33.955 137.255 34.125 ;
        RECT 137.545 33.955 137.715 34.125 ;
        RECT 138.005 33.955 138.175 34.125 ;
        RECT 138.465 33.955 138.635 34.125 ;
        RECT 138.925 33.955 139.095 34.125 ;
        RECT 139.385 33.955 139.555 34.125 ;
        RECT 139.845 33.955 140.015 34.125 ;
        RECT 140.305 33.955 140.475 34.125 ;
        RECT 140.765 33.955 140.935 34.125 ;
        RECT 141.225 33.955 141.395 34.125 ;
        RECT 141.685 33.955 141.855 34.125 ;
        RECT 142.145 33.955 142.315 34.125 ;
        RECT 142.605 33.955 142.775 34.125 ;
        RECT 143.065 33.955 143.235 34.125 ;
        RECT 143.525 33.955 143.695 34.125 ;
        RECT 143.985 33.955 144.155 34.125 ;
        RECT 55.665 28.515 55.835 28.685 ;
        RECT 56.125 28.515 56.295 28.685 ;
        RECT 56.585 28.515 56.755 28.685 ;
        RECT 57.045 28.515 57.215 28.685 ;
        RECT 57.505 28.515 57.675 28.685 ;
        RECT 57.965 28.515 58.135 28.685 ;
        RECT 58.425 28.515 58.595 28.685 ;
        RECT 58.885 28.515 59.055 28.685 ;
        RECT 59.345 28.515 59.515 28.685 ;
        RECT 59.805 28.515 59.975 28.685 ;
        RECT 60.265 28.515 60.435 28.685 ;
        RECT 60.725 28.515 60.895 28.685 ;
        RECT 61.185 28.515 61.355 28.685 ;
        RECT 61.645 28.515 61.815 28.685 ;
        RECT 62.105 28.515 62.275 28.685 ;
        RECT 62.565 28.515 62.735 28.685 ;
        RECT 63.025 28.515 63.195 28.685 ;
        RECT 63.485 28.515 63.655 28.685 ;
        RECT 63.945 28.515 64.115 28.685 ;
        RECT 64.405 28.515 64.575 28.685 ;
        RECT 64.865 28.515 65.035 28.685 ;
        RECT 65.325 28.515 65.495 28.685 ;
        RECT 65.785 28.515 65.955 28.685 ;
        RECT 66.245 28.515 66.415 28.685 ;
        RECT 66.705 28.515 66.875 28.685 ;
        RECT 67.165 28.515 67.335 28.685 ;
        RECT 67.625 28.515 67.795 28.685 ;
        RECT 68.085 28.515 68.255 28.685 ;
        RECT 68.545 28.515 68.715 28.685 ;
        RECT 69.005 28.515 69.175 28.685 ;
        RECT 69.465 28.515 69.635 28.685 ;
        RECT 69.925 28.515 70.095 28.685 ;
        RECT 70.385 28.515 70.555 28.685 ;
        RECT 70.845 28.515 71.015 28.685 ;
        RECT 71.305 28.515 71.475 28.685 ;
        RECT 71.765 28.515 71.935 28.685 ;
        RECT 72.225 28.515 72.395 28.685 ;
        RECT 72.685 28.515 72.855 28.685 ;
        RECT 73.145 28.515 73.315 28.685 ;
        RECT 73.605 28.515 73.775 28.685 ;
        RECT 74.065 28.515 74.235 28.685 ;
        RECT 74.525 28.515 74.695 28.685 ;
        RECT 74.985 28.515 75.155 28.685 ;
        RECT 75.445 28.515 75.615 28.685 ;
        RECT 75.905 28.515 76.075 28.685 ;
        RECT 76.365 28.515 76.535 28.685 ;
        RECT 76.825 28.515 76.995 28.685 ;
        RECT 77.285 28.515 77.455 28.685 ;
        RECT 77.745 28.515 77.915 28.685 ;
        RECT 78.205 28.515 78.375 28.685 ;
        RECT 78.665 28.515 78.835 28.685 ;
        RECT 79.125 28.515 79.295 28.685 ;
        RECT 79.585 28.515 79.755 28.685 ;
        RECT 80.045 28.515 80.215 28.685 ;
        RECT 80.505 28.515 80.675 28.685 ;
        RECT 80.965 28.515 81.135 28.685 ;
        RECT 81.425 28.515 81.595 28.685 ;
        RECT 81.885 28.515 82.055 28.685 ;
        RECT 82.345 28.515 82.515 28.685 ;
        RECT 82.805 28.515 82.975 28.685 ;
        RECT 83.265 28.515 83.435 28.685 ;
        RECT 83.725 28.515 83.895 28.685 ;
        RECT 84.185 28.515 84.355 28.685 ;
        RECT 84.645 28.515 84.815 28.685 ;
        RECT 85.105 28.515 85.275 28.685 ;
        RECT 85.565 28.515 85.735 28.685 ;
        RECT 86.025 28.515 86.195 28.685 ;
        RECT 86.485 28.515 86.655 28.685 ;
        RECT 86.945 28.515 87.115 28.685 ;
        RECT 87.405 28.515 87.575 28.685 ;
        RECT 87.865 28.515 88.035 28.685 ;
        RECT 88.325 28.515 88.495 28.685 ;
        RECT 88.785 28.515 88.955 28.685 ;
        RECT 89.245 28.515 89.415 28.685 ;
        RECT 89.705 28.515 89.875 28.685 ;
        RECT 90.165 28.515 90.335 28.685 ;
        RECT 90.625 28.515 90.795 28.685 ;
        RECT 91.085 28.515 91.255 28.685 ;
        RECT 91.545 28.515 91.715 28.685 ;
        RECT 92.005 28.515 92.175 28.685 ;
        RECT 92.465 28.515 92.635 28.685 ;
        RECT 92.925 28.515 93.095 28.685 ;
        RECT 93.385 28.515 93.555 28.685 ;
        RECT 93.845 28.515 94.015 28.685 ;
        RECT 94.305 28.515 94.475 28.685 ;
        RECT 94.765 28.515 94.935 28.685 ;
        RECT 95.225 28.515 95.395 28.685 ;
        RECT 95.685 28.515 95.855 28.685 ;
        RECT 96.145 28.515 96.315 28.685 ;
        RECT 96.605 28.515 96.775 28.685 ;
        RECT 97.065 28.515 97.235 28.685 ;
        RECT 97.525 28.515 97.695 28.685 ;
        RECT 97.985 28.515 98.155 28.685 ;
        RECT 98.445 28.515 98.615 28.685 ;
        RECT 98.905 28.515 99.075 28.685 ;
        RECT 99.365 28.515 99.535 28.685 ;
        RECT 99.825 28.515 99.995 28.685 ;
        RECT 100.285 28.515 100.455 28.685 ;
        RECT 100.745 28.515 100.915 28.685 ;
        RECT 101.205 28.515 101.375 28.685 ;
        RECT 101.665 28.515 101.835 28.685 ;
        RECT 102.125 28.515 102.295 28.685 ;
        RECT 102.585 28.515 102.755 28.685 ;
        RECT 103.045 28.515 103.215 28.685 ;
        RECT 103.505 28.515 103.675 28.685 ;
        RECT 103.965 28.515 104.135 28.685 ;
        RECT 104.425 28.515 104.595 28.685 ;
        RECT 104.885 28.515 105.055 28.685 ;
        RECT 105.345 28.515 105.515 28.685 ;
        RECT 105.805 28.515 105.975 28.685 ;
        RECT 106.265 28.515 106.435 28.685 ;
        RECT 106.725 28.515 106.895 28.685 ;
        RECT 107.185 28.515 107.355 28.685 ;
        RECT 107.645 28.515 107.815 28.685 ;
        RECT 108.105 28.515 108.275 28.685 ;
        RECT 108.565 28.515 108.735 28.685 ;
        RECT 109.025 28.515 109.195 28.685 ;
        RECT 109.485 28.515 109.655 28.685 ;
        RECT 109.945 28.515 110.115 28.685 ;
        RECT 110.405 28.515 110.575 28.685 ;
        RECT 110.865 28.515 111.035 28.685 ;
        RECT 111.325 28.515 111.495 28.685 ;
        RECT 111.785 28.515 111.955 28.685 ;
        RECT 112.245 28.515 112.415 28.685 ;
        RECT 112.705 28.515 112.875 28.685 ;
        RECT 113.165 28.515 113.335 28.685 ;
        RECT 113.625 28.515 113.795 28.685 ;
        RECT 114.085 28.515 114.255 28.685 ;
        RECT 114.545 28.515 114.715 28.685 ;
        RECT 115.005 28.515 115.175 28.685 ;
        RECT 115.465 28.515 115.635 28.685 ;
        RECT 115.925 28.515 116.095 28.685 ;
        RECT 116.385 28.515 116.555 28.685 ;
        RECT 116.845 28.515 117.015 28.685 ;
        RECT 117.305 28.515 117.475 28.685 ;
        RECT 117.765 28.515 117.935 28.685 ;
        RECT 118.225 28.515 118.395 28.685 ;
        RECT 118.685 28.515 118.855 28.685 ;
        RECT 119.145 28.515 119.315 28.685 ;
        RECT 119.605 28.515 119.775 28.685 ;
        RECT 120.065 28.515 120.235 28.685 ;
        RECT 120.525 28.515 120.695 28.685 ;
        RECT 120.985 28.515 121.155 28.685 ;
        RECT 121.445 28.515 121.615 28.685 ;
        RECT 121.905 28.515 122.075 28.685 ;
        RECT 122.365 28.515 122.535 28.685 ;
        RECT 122.825 28.515 122.995 28.685 ;
        RECT 123.285 28.515 123.455 28.685 ;
        RECT 123.745 28.515 123.915 28.685 ;
        RECT 124.205 28.515 124.375 28.685 ;
        RECT 124.665 28.515 124.835 28.685 ;
        RECT 125.125 28.515 125.295 28.685 ;
        RECT 125.585 28.515 125.755 28.685 ;
        RECT 126.045 28.515 126.215 28.685 ;
        RECT 126.505 28.515 126.675 28.685 ;
        RECT 126.965 28.515 127.135 28.685 ;
        RECT 127.425 28.515 127.595 28.685 ;
        RECT 127.885 28.515 128.055 28.685 ;
        RECT 128.345 28.515 128.515 28.685 ;
        RECT 128.805 28.515 128.975 28.685 ;
        RECT 129.265 28.515 129.435 28.685 ;
        RECT 129.725 28.515 129.895 28.685 ;
        RECT 130.185 28.515 130.355 28.685 ;
        RECT 130.645 28.515 130.815 28.685 ;
        RECT 131.105 28.515 131.275 28.685 ;
        RECT 131.565 28.515 131.735 28.685 ;
        RECT 132.025 28.515 132.195 28.685 ;
        RECT 132.485 28.515 132.655 28.685 ;
        RECT 132.945 28.515 133.115 28.685 ;
        RECT 133.405 28.515 133.575 28.685 ;
        RECT 133.865 28.515 134.035 28.685 ;
        RECT 134.325 28.515 134.495 28.685 ;
        RECT 134.785 28.515 134.955 28.685 ;
        RECT 135.245 28.515 135.415 28.685 ;
        RECT 135.705 28.515 135.875 28.685 ;
        RECT 136.165 28.515 136.335 28.685 ;
        RECT 136.625 28.515 136.795 28.685 ;
        RECT 137.085 28.515 137.255 28.685 ;
        RECT 137.545 28.515 137.715 28.685 ;
        RECT 138.005 28.515 138.175 28.685 ;
        RECT 138.465 28.515 138.635 28.685 ;
        RECT 138.925 28.515 139.095 28.685 ;
        RECT 139.385 28.515 139.555 28.685 ;
        RECT 139.845 28.515 140.015 28.685 ;
        RECT 140.305 28.515 140.475 28.685 ;
        RECT 140.765 28.515 140.935 28.685 ;
        RECT 141.225 28.515 141.395 28.685 ;
        RECT 141.685 28.515 141.855 28.685 ;
        RECT 142.145 28.515 142.315 28.685 ;
        RECT 142.605 28.515 142.775 28.685 ;
        RECT 143.065 28.515 143.235 28.685 ;
        RECT 143.525 28.515 143.695 28.685 ;
        RECT 143.985 28.515 144.155 28.685 ;
      LAYER met1 ;
        RECT 55.520 99.080 144.300 99.560 ;
        RECT 55.520 93.640 144.300 94.120 ;
        RECT 55.520 88.200 144.300 88.680 ;
        RECT 55.520 82.760 144.300 83.240 ;
        RECT 55.520 77.320 144.300 77.800 ;
        RECT 55.520 71.880 144.300 72.360 ;
        RECT 55.520 66.440 144.300 66.920 ;
        RECT 55.520 61.000 144.300 61.480 ;
        RECT 55.520 55.560 144.300 56.040 ;
        RECT 55.520 50.120 144.300 50.600 ;
        RECT 55.520 44.680 144.300 45.160 ;
        RECT 55.520 39.240 144.300 39.720 ;
        RECT 55.520 33.800 144.300 34.280 ;
        RECT 55.520 28.360 144.300 28.840 ;
      LAYER via ;
        RECT 65.845 99.190 66.105 99.450 ;
        RECT 66.165 99.190 66.425 99.450 ;
        RECT 66.485 99.190 66.745 99.450 ;
        RECT 66.805 99.190 67.065 99.450 ;
        RECT 67.125 99.190 67.385 99.450 ;
        RECT 88.040 99.190 88.300 99.450 ;
        RECT 88.360 99.190 88.620 99.450 ;
        RECT 88.680 99.190 88.940 99.450 ;
        RECT 89.000 99.190 89.260 99.450 ;
        RECT 89.320 99.190 89.580 99.450 ;
        RECT 110.235 99.190 110.495 99.450 ;
        RECT 110.555 99.190 110.815 99.450 ;
        RECT 110.875 99.190 111.135 99.450 ;
        RECT 111.195 99.190 111.455 99.450 ;
        RECT 111.515 99.190 111.775 99.450 ;
        RECT 132.430 99.190 132.690 99.450 ;
        RECT 132.750 99.190 133.010 99.450 ;
        RECT 133.070 99.190 133.330 99.450 ;
        RECT 133.390 99.190 133.650 99.450 ;
        RECT 133.710 99.190 133.970 99.450 ;
        RECT 65.845 93.750 66.105 94.010 ;
        RECT 66.165 93.750 66.425 94.010 ;
        RECT 66.485 93.750 66.745 94.010 ;
        RECT 66.805 93.750 67.065 94.010 ;
        RECT 67.125 93.750 67.385 94.010 ;
        RECT 88.040 93.750 88.300 94.010 ;
        RECT 88.360 93.750 88.620 94.010 ;
        RECT 88.680 93.750 88.940 94.010 ;
        RECT 89.000 93.750 89.260 94.010 ;
        RECT 89.320 93.750 89.580 94.010 ;
        RECT 110.235 93.750 110.495 94.010 ;
        RECT 110.555 93.750 110.815 94.010 ;
        RECT 110.875 93.750 111.135 94.010 ;
        RECT 111.195 93.750 111.455 94.010 ;
        RECT 111.515 93.750 111.775 94.010 ;
        RECT 132.430 93.750 132.690 94.010 ;
        RECT 132.750 93.750 133.010 94.010 ;
        RECT 133.070 93.750 133.330 94.010 ;
        RECT 133.390 93.750 133.650 94.010 ;
        RECT 133.710 93.750 133.970 94.010 ;
        RECT 65.845 88.310 66.105 88.570 ;
        RECT 66.165 88.310 66.425 88.570 ;
        RECT 66.485 88.310 66.745 88.570 ;
        RECT 66.805 88.310 67.065 88.570 ;
        RECT 67.125 88.310 67.385 88.570 ;
        RECT 88.040 88.310 88.300 88.570 ;
        RECT 88.360 88.310 88.620 88.570 ;
        RECT 88.680 88.310 88.940 88.570 ;
        RECT 89.000 88.310 89.260 88.570 ;
        RECT 89.320 88.310 89.580 88.570 ;
        RECT 110.235 88.310 110.495 88.570 ;
        RECT 110.555 88.310 110.815 88.570 ;
        RECT 110.875 88.310 111.135 88.570 ;
        RECT 111.195 88.310 111.455 88.570 ;
        RECT 111.515 88.310 111.775 88.570 ;
        RECT 132.430 88.310 132.690 88.570 ;
        RECT 132.750 88.310 133.010 88.570 ;
        RECT 133.070 88.310 133.330 88.570 ;
        RECT 133.390 88.310 133.650 88.570 ;
        RECT 133.710 88.310 133.970 88.570 ;
        RECT 65.845 82.870 66.105 83.130 ;
        RECT 66.165 82.870 66.425 83.130 ;
        RECT 66.485 82.870 66.745 83.130 ;
        RECT 66.805 82.870 67.065 83.130 ;
        RECT 67.125 82.870 67.385 83.130 ;
        RECT 88.040 82.870 88.300 83.130 ;
        RECT 88.360 82.870 88.620 83.130 ;
        RECT 88.680 82.870 88.940 83.130 ;
        RECT 89.000 82.870 89.260 83.130 ;
        RECT 89.320 82.870 89.580 83.130 ;
        RECT 110.235 82.870 110.495 83.130 ;
        RECT 110.555 82.870 110.815 83.130 ;
        RECT 110.875 82.870 111.135 83.130 ;
        RECT 111.195 82.870 111.455 83.130 ;
        RECT 111.515 82.870 111.775 83.130 ;
        RECT 132.430 82.870 132.690 83.130 ;
        RECT 132.750 82.870 133.010 83.130 ;
        RECT 133.070 82.870 133.330 83.130 ;
        RECT 133.390 82.870 133.650 83.130 ;
        RECT 133.710 82.870 133.970 83.130 ;
        RECT 65.845 77.430 66.105 77.690 ;
        RECT 66.165 77.430 66.425 77.690 ;
        RECT 66.485 77.430 66.745 77.690 ;
        RECT 66.805 77.430 67.065 77.690 ;
        RECT 67.125 77.430 67.385 77.690 ;
        RECT 88.040 77.430 88.300 77.690 ;
        RECT 88.360 77.430 88.620 77.690 ;
        RECT 88.680 77.430 88.940 77.690 ;
        RECT 89.000 77.430 89.260 77.690 ;
        RECT 89.320 77.430 89.580 77.690 ;
        RECT 110.235 77.430 110.495 77.690 ;
        RECT 110.555 77.430 110.815 77.690 ;
        RECT 110.875 77.430 111.135 77.690 ;
        RECT 111.195 77.430 111.455 77.690 ;
        RECT 111.515 77.430 111.775 77.690 ;
        RECT 132.430 77.430 132.690 77.690 ;
        RECT 132.750 77.430 133.010 77.690 ;
        RECT 133.070 77.430 133.330 77.690 ;
        RECT 133.390 77.430 133.650 77.690 ;
        RECT 133.710 77.430 133.970 77.690 ;
        RECT 65.845 71.990 66.105 72.250 ;
        RECT 66.165 71.990 66.425 72.250 ;
        RECT 66.485 71.990 66.745 72.250 ;
        RECT 66.805 71.990 67.065 72.250 ;
        RECT 67.125 71.990 67.385 72.250 ;
        RECT 88.040 71.990 88.300 72.250 ;
        RECT 88.360 71.990 88.620 72.250 ;
        RECT 88.680 71.990 88.940 72.250 ;
        RECT 89.000 71.990 89.260 72.250 ;
        RECT 89.320 71.990 89.580 72.250 ;
        RECT 110.235 71.990 110.495 72.250 ;
        RECT 110.555 71.990 110.815 72.250 ;
        RECT 110.875 71.990 111.135 72.250 ;
        RECT 111.195 71.990 111.455 72.250 ;
        RECT 111.515 71.990 111.775 72.250 ;
        RECT 132.430 71.990 132.690 72.250 ;
        RECT 132.750 71.990 133.010 72.250 ;
        RECT 133.070 71.990 133.330 72.250 ;
        RECT 133.390 71.990 133.650 72.250 ;
        RECT 133.710 71.990 133.970 72.250 ;
        RECT 65.845 66.550 66.105 66.810 ;
        RECT 66.165 66.550 66.425 66.810 ;
        RECT 66.485 66.550 66.745 66.810 ;
        RECT 66.805 66.550 67.065 66.810 ;
        RECT 67.125 66.550 67.385 66.810 ;
        RECT 88.040 66.550 88.300 66.810 ;
        RECT 88.360 66.550 88.620 66.810 ;
        RECT 88.680 66.550 88.940 66.810 ;
        RECT 89.000 66.550 89.260 66.810 ;
        RECT 89.320 66.550 89.580 66.810 ;
        RECT 110.235 66.550 110.495 66.810 ;
        RECT 110.555 66.550 110.815 66.810 ;
        RECT 110.875 66.550 111.135 66.810 ;
        RECT 111.195 66.550 111.455 66.810 ;
        RECT 111.515 66.550 111.775 66.810 ;
        RECT 132.430 66.550 132.690 66.810 ;
        RECT 132.750 66.550 133.010 66.810 ;
        RECT 133.070 66.550 133.330 66.810 ;
        RECT 133.390 66.550 133.650 66.810 ;
        RECT 133.710 66.550 133.970 66.810 ;
        RECT 65.845 61.110 66.105 61.370 ;
        RECT 66.165 61.110 66.425 61.370 ;
        RECT 66.485 61.110 66.745 61.370 ;
        RECT 66.805 61.110 67.065 61.370 ;
        RECT 67.125 61.110 67.385 61.370 ;
        RECT 88.040 61.110 88.300 61.370 ;
        RECT 88.360 61.110 88.620 61.370 ;
        RECT 88.680 61.110 88.940 61.370 ;
        RECT 89.000 61.110 89.260 61.370 ;
        RECT 89.320 61.110 89.580 61.370 ;
        RECT 110.235 61.110 110.495 61.370 ;
        RECT 110.555 61.110 110.815 61.370 ;
        RECT 110.875 61.110 111.135 61.370 ;
        RECT 111.195 61.110 111.455 61.370 ;
        RECT 111.515 61.110 111.775 61.370 ;
        RECT 132.430 61.110 132.690 61.370 ;
        RECT 132.750 61.110 133.010 61.370 ;
        RECT 133.070 61.110 133.330 61.370 ;
        RECT 133.390 61.110 133.650 61.370 ;
        RECT 133.710 61.110 133.970 61.370 ;
        RECT 65.845 55.670 66.105 55.930 ;
        RECT 66.165 55.670 66.425 55.930 ;
        RECT 66.485 55.670 66.745 55.930 ;
        RECT 66.805 55.670 67.065 55.930 ;
        RECT 67.125 55.670 67.385 55.930 ;
        RECT 88.040 55.670 88.300 55.930 ;
        RECT 88.360 55.670 88.620 55.930 ;
        RECT 88.680 55.670 88.940 55.930 ;
        RECT 89.000 55.670 89.260 55.930 ;
        RECT 89.320 55.670 89.580 55.930 ;
        RECT 110.235 55.670 110.495 55.930 ;
        RECT 110.555 55.670 110.815 55.930 ;
        RECT 110.875 55.670 111.135 55.930 ;
        RECT 111.195 55.670 111.455 55.930 ;
        RECT 111.515 55.670 111.775 55.930 ;
        RECT 132.430 55.670 132.690 55.930 ;
        RECT 132.750 55.670 133.010 55.930 ;
        RECT 133.070 55.670 133.330 55.930 ;
        RECT 133.390 55.670 133.650 55.930 ;
        RECT 133.710 55.670 133.970 55.930 ;
        RECT 65.845 50.230 66.105 50.490 ;
        RECT 66.165 50.230 66.425 50.490 ;
        RECT 66.485 50.230 66.745 50.490 ;
        RECT 66.805 50.230 67.065 50.490 ;
        RECT 67.125 50.230 67.385 50.490 ;
        RECT 88.040 50.230 88.300 50.490 ;
        RECT 88.360 50.230 88.620 50.490 ;
        RECT 88.680 50.230 88.940 50.490 ;
        RECT 89.000 50.230 89.260 50.490 ;
        RECT 89.320 50.230 89.580 50.490 ;
        RECT 110.235 50.230 110.495 50.490 ;
        RECT 110.555 50.230 110.815 50.490 ;
        RECT 110.875 50.230 111.135 50.490 ;
        RECT 111.195 50.230 111.455 50.490 ;
        RECT 111.515 50.230 111.775 50.490 ;
        RECT 132.430 50.230 132.690 50.490 ;
        RECT 132.750 50.230 133.010 50.490 ;
        RECT 133.070 50.230 133.330 50.490 ;
        RECT 133.390 50.230 133.650 50.490 ;
        RECT 133.710 50.230 133.970 50.490 ;
        RECT 65.845 44.790 66.105 45.050 ;
        RECT 66.165 44.790 66.425 45.050 ;
        RECT 66.485 44.790 66.745 45.050 ;
        RECT 66.805 44.790 67.065 45.050 ;
        RECT 67.125 44.790 67.385 45.050 ;
        RECT 88.040 44.790 88.300 45.050 ;
        RECT 88.360 44.790 88.620 45.050 ;
        RECT 88.680 44.790 88.940 45.050 ;
        RECT 89.000 44.790 89.260 45.050 ;
        RECT 89.320 44.790 89.580 45.050 ;
        RECT 110.235 44.790 110.495 45.050 ;
        RECT 110.555 44.790 110.815 45.050 ;
        RECT 110.875 44.790 111.135 45.050 ;
        RECT 111.195 44.790 111.455 45.050 ;
        RECT 111.515 44.790 111.775 45.050 ;
        RECT 132.430 44.790 132.690 45.050 ;
        RECT 132.750 44.790 133.010 45.050 ;
        RECT 133.070 44.790 133.330 45.050 ;
        RECT 133.390 44.790 133.650 45.050 ;
        RECT 133.710 44.790 133.970 45.050 ;
        RECT 65.845 39.350 66.105 39.610 ;
        RECT 66.165 39.350 66.425 39.610 ;
        RECT 66.485 39.350 66.745 39.610 ;
        RECT 66.805 39.350 67.065 39.610 ;
        RECT 67.125 39.350 67.385 39.610 ;
        RECT 88.040 39.350 88.300 39.610 ;
        RECT 88.360 39.350 88.620 39.610 ;
        RECT 88.680 39.350 88.940 39.610 ;
        RECT 89.000 39.350 89.260 39.610 ;
        RECT 89.320 39.350 89.580 39.610 ;
        RECT 110.235 39.350 110.495 39.610 ;
        RECT 110.555 39.350 110.815 39.610 ;
        RECT 110.875 39.350 111.135 39.610 ;
        RECT 111.195 39.350 111.455 39.610 ;
        RECT 111.515 39.350 111.775 39.610 ;
        RECT 132.430 39.350 132.690 39.610 ;
        RECT 132.750 39.350 133.010 39.610 ;
        RECT 133.070 39.350 133.330 39.610 ;
        RECT 133.390 39.350 133.650 39.610 ;
        RECT 133.710 39.350 133.970 39.610 ;
        RECT 65.845 33.910 66.105 34.170 ;
        RECT 66.165 33.910 66.425 34.170 ;
        RECT 66.485 33.910 66.745 34.170 ;
        RECT 66.805 33.910 67.065 34.170 ;
        RECT 67.125 33.910 67.385 34.170 ;
        RECT 88.040 33.910 88.300 34.170 ;
        RECT 88.360 33.910 88.620 34.170 ;
        RECT 88.680 33.910 88.940 34.170 ;
        RECT 89.000 33.910 89.260 34.170 ;
        RECT 89.320 33.910 89.580 34.170 ;
        RECT 110.235 33.910 110.495 34.170 ;
        RECT 110.555 33.910 110.815 34.170 ;
        RECT 110.875 33.910 111.135 34.170 ;
        RECT 111.195 33.910 111.455 34.170 ;
        RECT 111.515 33.910 111.775 34.170 ;
        RECT 132.430 33.910 132.690 34.170 ;
        RECT 132.750 33.910 133.010 34.170 ;
        RECT 133.070 33.910 133.330 34.170 ;
        RECT 133.390 33.910 133.650 34.170 ;
        RECT 133.710 33.910 133.970 34.170 ;
        RECT 65.845 28.470 66.105 28.730 ;
        RECT 66.165 28.470 66.425 28.730 ;
        RECT 66.485 28.470 66.745 28.730 ;
        RECT 66.805 28.470 67.065 28.730 ;
        RECT 67.125 28.470 67.385 28.730 ;
        RECT 88.040 28.470 88.300 28.730 ;
        RECT 88.360 28.470 88.620 28.730 ;
        RECT 88.680 28.470 88.940 28.730 ;
        RECT 89.000 28.470 89.260 28.730 ;
        RECT 89.320 28.470 89.580 28.730 ;
        RECT 110.235 28.470 110.495 28.730 ;
        RECT 110.555 28.470 110.815 28.730 ;
        RECT 110.875 28.470 111.135 28.730 ;
        RECT 111.195 28.470 111.455 28.730 ;
        RECT 111.515 28.470 111.775 28.730 ;
        RECT 132.430 28.470 132.690 28.730 ;
        RECT 132.750 28.470 133.010 28.730 ;
        RECT 133.070 28.470 133.330 28.730 ;
        RECT 133.390 28.470 133.650 28.730 ;
        RECT 133.710 28.470 133.970 28.730 ;
      LAYER met2 ;
        RECT 65.845 99.135 67.385 99.505 ;
        RECT 88.040 99.135 89.580 99.505 ;
        RECT 110.235 99.135 111.775 99.505 ;
        RECT 132.430 99.135 133.970 99.505 ;
        RECT 65.845 93.695 67.385 94.065 ;
        RECT 88.040 93.695 89.580 94.065 ;
        RECT 110.235 93.695 111.775 94.065 ;
        RECT 132.430 93.695 133.970 94.065 ;
        RECT 65.845 88.255 67.385 88.625 ;
        RECT 88.040 88.255 89.580 88.625 ;
        RECT 110.235 88.255 111.775 88.625 ;
        RECT 132.430 88.255 133.970 88.625 ;
        RECT 65.845 82.815 67.385 83.185 ;
        RECT 88.040 82.815 89.580 83.185 ;
        RECT 110.235 82.815 111.775 83.185 ;
        RECT 132.430 82.815 133.970 83.185 ;
        RECT 65.845 77.375 67.385 77.745 ;
        RECT 88.040 77.375 89.580 77.745 ;
        RECT 110.235 77.375 111.775 77.745 ;
        RECT 132.430 77.375 133.970 77.745 ;
        RECT 65.845 71.935 67.385 72.305 ;
        RECT 88.040 71.935 89.580 72.305 ;
        RECT 110.235 71.935 111.775 72.305 ;
        RECT 132.430 71.935 133.970 72.305 ;
        RECT 65.845 66.495 67.385 66.865 ;
        RECT 88.040 66.495 89.580 66.865 ;
        RECT 110.235 66.495 111.775 66.865 ;
        RECT 132.430 66.495 133.970 66.865 ;
        RECT 65.845 61.055 67.385 61.425 ;
        RECT 88.040 61.055 89.580 61.425 ;
        RECT 110.235 61.055 111.775 61.425 ;
        RECT 132.430 61.055 133.970 61.425 ;
        RECT 65.845 55.615 67.385 55.985 ;
        RECT 88.040 55.615 89.580 55.985 ;
        RECT 110.235 55.615 111.775 55.985 ;
        RECT 132.430 55.615 133.970 55.985 ;
        RECT 65.845 50.175 67.385 50.545 ;
        RECT 88.040 50.175 89.580 50.545 ;
        RECT 110.235 50.175 111.775 50.545 ;
        RECT 132.430 50.175 133.970 50.545 ;
        RECT 65.845 44.735 67.385 45.105 ;
        RECT 88.040 44.735 89.580 45.105 ;
        RECT 110.235 44.735 111.775 45.105 ;
        RECT 132.430 44.735 133.970 45.105 ;
        RECT 65.845 39.295 67.385 39.665 ;
        RECT 88.040 39.295 89.580 39.665 ;
        RECT 110.235 39.295 111.775 39.665 ;
        RECT 132.430 39.295 133.970 39.665 ;
        RECT 65.845 33.855 67.385 34.225 ;
        RECT 88.040 33.855 89.580 34.225 ;
        RECT 110.235 33.855 111.775 34.225 ;
        RECT 132.430 33.855 133.970 34.225 ;
        RECT 65.845 28.415 67.385 28.785 ;
        RECT 88.040 28.415 89.580 28.785 ;
        RECT 110.235 28.415 111.775 28.785 ;
        RECT 132.430 28.415 133.970 28.785 ;
      LAYER via2 ;
        RECT 65.875 99.180 66.155 99.460 ;
        RECT 66.275 99.180 66.555 99.460 ;
        RECT 66.675 99.180 66.955 99.460 ;
        RECT 67.075 99.180 67.355 99.460 ;
        RECT 88.070 99.180 88.350 99.460 ;
        RECT 88.470 99.180 88.750 99.460 ;
        RECT 88.870 99.180 89.150 99.460 ;
        RECT 89.270 99.180 89.550 99.460 ;
        RECT 110.265 99.180 110.545 99.460 ;
        RECT 110.665 99.180 110.945 99.460 ;
        RECT 111.065 99.180 111.345 99.460 ;
        RECT 111.465 99.180 111.745 99.460 ;
        RECT 132.460 99.180 132.740 99.460 ;
        RECT 132.860 99.180 133.140 99.460 ;
        RECT 133.260 99.180 133.540 99.460 ;
        RECT 133.660 99.180 133.940 99.460 ;
        RECT 65.875 93.740 66.155 94.020 ;
        RECT 66.275 93.740 66.555 94.020 ;
        RECT 66.675 93.740 66.955 94.020 ;
        RECT 67.075 93.740 67.355 94.020 ;
        RECT 88.070 93.740 88.350 94.020 ;
        RECT 88.470 93.740 88.750 94.020 ;
        RECT 88.870 93.740 89.150 94.020 ;
        RECT 89.270 93.740 89.550 94.020 ;
        RECT 110.265 93.740 110.545 94.020 ;
        RECT 110.665 93.740 110.945 94.020 ;
        RECT 111.065 93.740 111.345 94.020 ;
        RECT 111.465 93.740 111.745 94.020 ;
        RECT 132.460 93.740 132.740 94.020 ;
        RECT 132.860 93.740 133.140 94.020 ;
        RECT 133.260 93.740 133.540 94.020 ;
        RECT 133.660 93.740 133.940 94.020 ;
        RECT 65.875 88.300 66.155 88.580 ;
        RECT 66.275 88.300 66.555 88.580 ;
        RECT 66.675 88.300 66.955 88.580 ;
        RECT 67.075 88.300 67.355 88.580 ;
        RECT 88.070 88.300 88.350 88.580 ;
        RECT 88.470 88.300 88.750 88.580 ;
        RECT 88.870 88.300 89.150 88.580 ;
        RECT 89.270 88.300 89.550 88.580 ;
        RECT 110.265 88.300 110.545 88.580 ;
        RECT 110.665 88.300 110.945 88.580 ;
        RECT 111.065 88.300 111.345 88.580 ;
        RECT 111.465 88.300 111.745 88.580 ;
        RECT 132.460 88.300 132.740 88.580 ;
        RECT 132.860 88.300 133.140 88.580 ;
        RECT 133.260 88.300 133.540 88.580 ;
        RECT 133.660 88.300 133.940 88.580 ;
        RECT 65.875 82.860 66.155 83.140 ;
        RECT 66.275 82.860 66.555 83.140 ;
        RECT 66.675 82.860 66.955 83.140 ;
        RECT 67.075 82.860 67.355 83.140 ;
        RECT 88.070 82.860 88.350 83.140 ;
        RECT 88.470 82.860 88.750 83.140 ;
        RECT 88.870 82.860 89.150 83.140 ;
        RECT 89.270 82.860 89.550 83.140 ;
        RECT 110.265 82.860 110.545 83.140 ;
        RECT 110.665 82.860 110.945 83.140 ;
        RECT 111.065 82.860 111.345 83.140 ;
        RECT 111.465 82.860 111.745 83.140 ;
        RECT 132.460 82.860 132.740 83.140 ;
        RECT 132.860 82.860 133.140 83.140 ;
        RECT 133.260 82.860 133.540 83.140 ;
        RECT 133.660 82.860 133.940 83.140 ;
        RECT 65.875 77.420 66.155 77.700 ;
        RECT 66.275 77.420 66.555 77.700 ;
        RECT 66.675 77.420 66.955 77.700 ;
        RECT 67.075 77.420 67.355 77.700 ;
        RECT 88.070 77.420 88.350 77.700 ;
        RECT 88.470 77.420 88.750 77.700 ;
        RECT 88.870 77.420 89.150 77.700 ;
        RECT 89.270 77.420 89.550 77.700 ;
        RECT 110.265 77.420 110.545 77.700 ;
        RECT 110.665 77.420 110.945 77.700 ;
        RECT 111.065 77.420 111.345 77.700 ;
        RECT 111.465 77.420 111.745 77.700 ;
        RECT 132.460 77.420 132.740 77.700 ;
        RECT 132.860 77.420 133.140 77.700 ;
        RECT 133.260 77.420 133.540 77.700 ;
        RECT 133.660 77.420 133.940 77.700 ;
        RECT 65.875 71.980 66.155 72.260 ;
        RECT 66.275 71.980 66.555 72.260 ;
        RECT 66.675 71.980 66.955 72.260 ;
        RECT 67.075 71.980 67.355 72.260 ;
        RECT 88.070 71.980 88.350 72.260 ;
        RECT 88.470 71.980 88.750 72.260 ;
        RECT 88.870 71.980 89.150 72.260 ;
        RECT 89.270 71.980 89.550 72.260 ;
        RECT 110.265 71.980 110.545 72.260 ;
        RECT 110.665 71.980 110.945 72.260 ;
        RECT 111.065 71.980 111.345 72.260 ;
        RECT 111.465 71.980 111.745 72.260 ;
        RECT 132.460 71.980 132.740 72.260 ;
        RECT 132.860 71.980 133.140 72.260 ;
        RECT 133.260 71.980 133.540 72.260 ;
        RECT 133.660 71.980 133.940 72.260 ;
        RECT 65.875 66.540 66.155 66.820 ;
        RECT 66.275 66.540 66.555 66.820 ;
        RECT 66.675 66.540 66.955 66.820 ;
        RECT 67.075 66.540 67.355 66.820 ;
        RECT 88.070 66.540 88.350 66.820 ;
        RECT 88.470 66.540 88.750 66.820 ;
        RECT 88.870 66.540 89.150 66.820 ;
        RECT 89.270 66.540 89.550 66.820 ;
        RECT 110.265 66.540 110.545 66.820 ;
        RECT 110.665 66.540 110.945 66.820 ;
        RECT 111.065 66.540 111.345 66.820 ;
        RECT 111.465 66.540 111.745 66.820 ;
        RECT 132.460 66.540 132.740 66.820 ;
        RECT 132.860 66.540 133.140 66.820 ;
        RECT 133.260 66.540 133.540 66.820 ;
        RECT 133.660 66.540 133.940 66.820 ;
        RECT 65.875 61.100 66.155 61.380 ;
        RECT 66.275 61.100 66.555 61.380 ;
        RECT 66.675 61.100 66.955 61.380 ;
        RECT 67.075 61.100 67.355 61.380 ;
        RECT 88.070 61.100 88.350 61.380 ;
        RECT 88.470 61.100 88.750 61.380 ;
        RECT 88.870 61.100 89.150 61.380 ;
        RECT 89.270 61.100 89.550 61.380 ;
        RECT 110.265 61.100 110.545 61.380 ;
        RECT 110.665 61.100 110.945 61.380 ;
        RECT 111.065 61.100 111.345 61.380 ;
        RECT 111.465 61.100 111.745 61.380 ;
        RECT 132.460 61.100 132.740 61.380 ;
        RECT 132.860 61.100 133.140 61.380 ;
        RECT 133.260 61.100 133.540 61.380 ;
        RECT 133.660 61.100 133.940 61.380 ;
        RECT 65.875 55.660 66.155 55.940 ;
        RECT 66.275 55.660 66.555 55.940 ;
        RECT 66.675 55.660 66.955 55.940 ;
        RECT 67.075 55.660 67.355 55.940 ;
        RECT 88.070 55.660 88.350 55.940 ;
        RECT 88.470 55.660 88.750 55.940 ;
        RECT 88.870 55.660 89.150 55.940 ;
        RECT 89.270 55.660 89.550 55.940 ;
        RECT 110.265 55.660 110.545 55.940 ;
        RECT 110.665 55.660 110.945 55.940 ;
        RECT 111.065 55.660 111.345 55.940 ;
        RECT 111.465 55.660 111.745 55.940 ;
        RECT 132.460 55.660 132.740 55.940 ;
        RECT 132.860 55.660 133.140 55.940 ;
        RECT 133.260 55.660 133.540 55.940 ;
        RECT 133.660 55.660 133.940 55.940 ;
        RECT 65.875 50.220 66.155 50.500 ;
        RECT 66.275 50.220 66.555 50.500 ;
        RECT 66.675 50.220 66.955 50.500 ;
        RECT 67.075 50.220 67.355 50.500 ;
        RECT 88.070 50.220 88.350 50.500 ;
        RECT 88.470 50.220 88.750 50.500 ;
        RECT 88.870 50.220 89.150 50.500 ;
        RECT 89.270 50.220 89.550 50.500 ;
        RECT 110.265 50.220 110.545 50.500 ;
        RECT 110.665 50.220 110.945 50.500 ;
        RECT 111.065 50.220 111.345 50.500 ;
        RECT 111.465 50.220 111.745 50.500 ;
        RECT 132.460 50.220 132.740 50.500 ;
        RECT 132.860 50.220 133.140 50.500 ;
        RECT 133.260 50.220 133.540 50.500 ;
        RECT 133.660 50.220 133.940 50.500 ;
        RECT 65.875 44.780 66.155 45.060 ;
        RECT 66.275 44.780 66.555 45.060 ;
        RECT 66.675 44.780 66.955 45.060 ;
        RECT 67.075 44.780 67.355 45.060 ;
        RECT 88.070 44.780 88.350 45.060 ;
        RECT 88.470 44.780 88.750 45.060 ;
        RECT 88.870 44.780 89.150 45.060 ;
        RECT 89.270 44.780 89.550 45.060 ;
        RECT 110.265 44.780 110.545 45.060 ;
        RECT 110.665 44.780 110.945 45.060 ;
        RECT 111.065 44.780 111.345 45.060 ;
        RECT 111.465 44.780 111.745 45.060 ;
        RECT 132.460 44.780 132.740 45.060 ;
        RECT 132.860 44.780 133.140 45.060 ;
        RECT 133.260 44.780 133.540 45.060 ;
        RECT 133.660 44.780 133.940 45.060 ;
        RECT 65.875 39.340 66.155 39.620 ;
        RECT 66.275 39.340 66.555 39.620 ;
        RECT 66.675 39.340 66.955 39.620 ;
        RECT 67.075 39.340 67.355 39.620 ;
        RECT 88.070 39.340 88.350 39.620 ;
        RECT 88.470 39.340 88.750 39.620 ;
        RECT 88.870 39.340 89.150 39.620 ;
        RECT 89.270 39.340 89.550 39.620 ;
        RECT 110.265 39.340 110.545 39.620 ;
        RECT 110.665 39.340 110.945 39.620 ;
        RECT 111.065 39.340 111.345 39.620 ;
        RECT 111.465 39.340 111.745 39.620 ;
        RECT 132.460 39.340 132.740 39.620 ;
        RECT 132.860 39.340 133.140 39.620 ;
        RECT 133.260 39.340 133.540 39.620 ;
        RECT 133.660 39.340 133.940 39.620 ;
        RECT 65.875 33.900 66.155 34.180 ;
        RECT 66.275 33.900 66.555 34.180 ;
        RECT 66.675 33.900 66.955 34.180 ;
        RECT 67.075 33.900 67.355 34.180 ;
        RECT 88.070 33.900 88.350 34.180 ;
        RECT 88.470 33.900 88.750 34.180 ;
        RECT 88.870 33.900 89.150 34.180 ;
        RECT 89.270 33.900 89.550 34.180 ;
        RECT 110.265 33.900 110.545 34.180 ;
        RECT 110.665 33.900 110.945 34.180 ;
        RECT 111.065 33.900 111.345 34.180 ;
        RECT 111.465 33.900 111.745 34.180 ;
        RECT 132.460 33.900 132.740 34.180 ;
        RECT 132.860 33.900 133.140 34.180 ;
        RECT 133.260 33.900 133.540 34.180 ;
        RECT 133.660 33.900 133.940 34.180 ;
        RECT 65.875 28.460 66.155 28.740 ;
        RECT 66.275 28.460 66.555 28.740 ;
        RECT 66.675 28.460 66.955 28.740 ;
        RECT 67.075 28.460 67.355 28.740 ;
        RECT 88.070 28.460 88.350 28.740 ;
        RECT 88.470 28.460 88.750 28.740 ;
        RECT 88.870 28.460 89.150 28.740 ;
        RECT 89.270 28.460 89.550 28.740 ;
        RECT 110.265 28.460 110.545 28.740 ;
        RECT 110.665 28.460 110.945 28.740 ;
        RECT 111.065 28.460 111.345 28.740 ;
        RECT 111.465 28.460 111.745 28.740 ;
        RECT 132.460 28.460 132.740 28.740 ;
        RECT 132.860 28.460 133.140 28.740 ;
        RECT 133.260 28.460 133.540 28.740 ;
        RECT 133.660 28.460 133.940 28.740 ;
      LAYER met3 ;
        RECT 65.825 99.155 67.405 99.485 ;
        RECT 88.020 99.155 89.600 99.485 ;
        RECT 110.215 99.155 111.795 99.485 ;
        RECT 132.410 99.155 133.990 99.485 ;
        RECT 65.825 93.715 67.405 94.045 ;
        RECT 88.020 93.715 89.600 94.045 ;
        RECT 110.215 93.715 111.795 94.045 ;
        RECT 132.410 93.715 133.990 94.045 ;
        RECT 65.825 88.275 67.405 88.605 ;
        RECT 88.020 88.275 89.600 88.605 ;
        RECT 110.215 88.275 111.795 88.605 ;
        RECT 132.410 88.275 133.990 88.605 ;
        RECT 65.825 82.835 67.405 83.165 ;
        RECT 88.020 82.835 89.600 83.165 ;
        RECT 110.215 82.835 111.795 83.165 ;
        RECT 132.410 82.835 133.990 83.165 ;
        RECT 65.825 77.395 67.405 77.725 ;
        RECT 88.020 77.395 89.600 77.725 ;
        RECT 110.215 77.395 111.795 77.725 ;
        RECT 132.410 77.395 133.990 77.725 ;
        RECT 65.825 71.955 67.405 72.285 ;
        RECT 88.020 71.955 89.600 72.285 ;
        RECT 110.215 71.955 111.795 72.285 ;
        RECT 132.410 71.955 133.990 72.285 ;
        RECT 65.825 66.515 67.405 66.845 ;
        RECT 88.020 66.515 89.600 66.845 ;
        RECT 110.215 66.515 111.795 66.845 ;
        RECT 132.410 66.515 133.990 66.845 ;
        RECT 65.825 61.075 67.405 61.405 ;
        RECT 88.020 61.075 89.600 61.405 ;
        RECT 110.215 61.075 111.795 61.405 ;
        RECT 132.410 61.075 133.990 61.405 ;
        RECT 65.825 55.635 67.405 55.965 ;
        RECT 88.020 55.635 89.600 55.965 ;
        RECT 110.215 55.635 111.795 55.965 ;
        RECT 132.410 55.635 133.990 55.965 ;
        RECT 65.825 50.195 67.405 50.525 ;
        RECT 88.020 50.195 89.600 50.525 ;
        RECT 110.215 50.195 111.795 50.525 ;
        RECT 132.410 50.195 133.990 50.525 ;
        RECT 65.825 44.755 67.405 45.085 ;
        RECT 88.020 44.755 89.600 45.085 ;
        RECT 110.215 44.755 111.795 45.085 ;
        RECT 132.410 44.755 133.990 45.085 ;
        RECT 65.825 39.315 67.405 39.645 ;
        RECT 88.020 39.315 89.600 39.645 ;
        RECT 110.215 39.315 111.795 39.645 ;
        RECT 132.410 39.315 133.990 39.645 ;
        RECT 65.825 33.875 67.405 34.205 ;
        RECT 88.020 33.875 89.600 34.205 ;
        RECT 110.215 33.875 111.795 34.205 ;
        RECT 132.410 33.875 133.990 34.205 ;
        RECT 65.825 28.435 67.405 28.765 ;
        RECT 88.020 28.435 89.600 28.765 ;
        RECT 110.215 28.435 111.795 28.765 ;
        RECT 132.410 28.435 133.990 28.765 ;
      LAYER via3 ;
        RECT 65.855 99.160 66.175 99.480 ;
        RECT 66.255 99.160 66.575 99.480 ;
        RECT 66.655 99.160 66.975 99.480 ;
        RECT 67.055 99.160 67.375 99.480 ;
        RECT 88.050 99.160 88.370 99.480 ;
        RECT 88.450 99.160 88.770 99.480 ;
        RECT 88.850 99.160 89.170 99.480 ;
        RECT 89.250 99.160 89.570 99.480 ;
        RECT 110.245 99.160 110.565 99.480 ;
        RECT 110.645 99.160 110.965 99.480 ;
        RECT 111.045 99.160 111.365 99.480 ;
        RECT 111.445 99.160 111.765 99.480 ;
        RECT 132.440 99.160 132.760 99.480 ;
        RECT 132.840 99.160 133.160 99.480 ;
        RECT 133.240 99.160 133.560 99.480 ;
        RECT 133.640 99.160 133.960 99.480 ;
        RECT 65.855 93.720 66.175 94.040 ;
        RECT 66.255 93.720 66.575 94.040 ;
        RECT 66.655 93.720 66.975 94.040 ;
        RECT 67.055 93.720 67.375 94.040 ;
        RECT 88.050 93.720 88.370 94.040 ;
        RECT 88.450 93.720 88.770 94.040 ;
        RECT 88.850 93.720 89.170 94.040 ;
        RECT 89.250 93.720 89.570 94.040 ;
        RECT 110.245 93.720 110.565 94.040 ;
        RECT 110.645 93.720 110.965 94.040 ;
        RECT 111.045 93.720 111.365 94.040 ;
        RECT 111.445 93.720 111.765 94.040 ;
        RECT 132.440 93.720 132.760 94.040 ;
        RECT 132.840 93.720 133.160 94.040 ;
        RECT 133.240 93.720 133.560 94.040 ;
        RECT 133.640 93.720 133.960 94.040 ;
        RECT 65.855 88.280 66.175 88.600 ;
        RECT 66.255 88.280 66.575 88.600 ;
        RECT 66.655 88.280 66.975 88.600 ;
        RECT 67.055 88.280 67.375 88.600 ;
        RECT 88.050 88.280 88.370 88.600 ;
        RECT 88.450 88.280 88.770 88.600 ;
        RECT 88.850 88.280 89.170 88.600 ;
        RECT 89.250 88.280 89.570 88.600 ;
        RECT 110.245 88.280 110.565 88.600 ;
        RECT 110.645 88.280 110.965 88.600 ;
        RECT 111.045 88.280 111.365 88.600 ;
        RECT 111.445 88.280 111.765 88.600 ;
        RECT 132.440 88.280 132.760 88.600 ;
        RECT 132.840 88.280 133.160 88.600 ;
        RECT 133.240 88.280 133.560 88.600 ;
        RECT 133.640 88.280 133.960 88.600 ;
        RECT 65.855 82.840 66.175 83.160 ;
        RECT 66.255 82.840 66.575 83.160 ;
        RECT 66.655 82.840 66.975 83.160 ;
        RECT 67.055 82.840 67.375 83.160 ;
        RECT 88.050 82.840 88.370 83.160 ;
        RECT 88.450 82.840 88.770 83.160 ;
        RECT 88.850 82.840 89.170 83.160 ;
        RECT 89.250 82.840 89.570 83.160 ;
        RECT 110.245 82.840 110.565 83.160 ;
        RECT 110.645 82.840 110.965 83.160 ;
        RECT 111.045 82.840 111.365 83.160 ;
        RECT 111.445 82.840 111.765 83.160 ;
        RECT 132.440 82.840 132.760 83.160 ;
        RECT 132.840 82.840 133.160 83.160 ;
        RECT 133.240 82.840 133.560 83.160 ;
        RECT 133.640 82.840 133.960 83.160 ;
        RECT 65.855 77.400 66.175 77.720 ;
        RECT 66.255 77.400 66.575 77.720 ;
        RECT 66.655 77.400 66.975 77.720 ;
        RECT 67.055 77.400 67.375 77.720 ;
        RECT 88.050 77.400 88.370 77.720 ;
        RECT 88.450 77.400 88.770 77.720 ;
        RECT 88.850 77.400 89.170 77.720 ;
        RECT 89.250 77.400 89.570 77.720 ;
        RECT 110.245 77.400 110.565 77.720 ;
        RECT 110.645 77.400 110.965 77.720 ;
        RECT 111.045 77.400 111.365 77.720 ;
        RECT 111.445 77.400 111.765 77.720 ;
        RECT 132.440 77.400 132.760 77.720 ;
        RECT 132.840 77.400 133.160 77.720 ;
        RECT 133.240 77.400 133.560 77.720 ;
        RECT 133.640 77.400 133.960 77.720 ;
        RECT 65.855 71.960 66.175 72.280 ;
        RECT 66.255 71.960 66.575 72.280 ;
        RECT 66.655 71.960 66.975 72.280 ;
        RECT 67.055 71.960 67.375 72.280 ;
        RECT 88.050 71.960 88.370 72.280 ;
        RECT 88.450 71.960 88.770 72.280 ;
        RECT 88.850 71.960 89.170 72.280 ;
        RECT 89.250 71.960 89.570 72.280 ;
        RECT 110.245 71.960 110.565 72.280 ;
        RECT 110.645 71.960 110.965 72.280 ;
        RECT 111.045 71.960 111.365 72.280 ;
        RECT 111.445 71.960 111.765 72.280 ;
        RECT 132.440 71.960 132.760 72.280 ;
        RECT 132.840 71.960 133.160 72.280 ;
        RECT 133.240 71.960 133.560 72.280 ;
        RECT 133.640 71.960 133.960 72.280 ;
        RECT 65.855 66.520 66.175 66.840 ;
        RECT 66.255 66.520 66.575 66.840 ;
        RECT 66.655 66.520 66.975 66.840 ;
        RECT 67.055 66.520 67.375 66.840 ;
        RECT 88.050 66.520 88.370 66.840 ;
        RECT 88.450 66.520 88.770 66.840 ;
        RECT 88.850 66.520 89.170 66.840 ;
        RECT 89.250 66.520 89.570 66.840 ;
        RECT 110.245 66.520 110.565 66.840 ;
        RECT 110.645 66.520 110.965 66.840 ;
        RECT 111.045 66.520 111.365 66.840 ;
        RECT 111.445 66.520 111.765 66.840 ;
        RECT 132.440 66.520 132.760 66.840 ;
        RECT 132.840 66.520 133.160 66.840 ;
        RECT 133.240 66.520 133.560 66.840 ;
        RECT 133.640 66.520 133.960 66.840 ;
        RECT 65.855 61.080 66.175 61.400 ;
        RECT 66.255 61.080 66.575 61.400 ;
        RECT 66.655 61.080 66.975 61.400 ;
        RECT 67.055 61.080 67.375 61.400 ;
        RECT 88.050 61.080 88.370 61.400 ;
        RECT 88.450 61.080 88.770 61.400 ;
        RECT 88.850 61.080 89.170 61.400 ;
        RECT 89.250 61.080 89.570 61.400 ;
        RECT 110.245 61.080 110.565 61.400 ;
        RECT 110.645 61.080 110.965 61.400 ;
        RECT 111.045 61.080 111.365 61.400 ;
        RECT 111.445 61.080 111.765 61.400 ;
        RECT 132.440 61.080 132.760 61.400 ;
        RECT 132.840 61.080 133.160 61.400 ;
        RECT 133.240 61.080 133.560 61.400 ;
        RECT 133.640 61.080 133.960 61.400 ;
        RECT 65.855 55.640 66.175 55.960 ;
        RECT 66.255 55.640 66.575 55.960 ;
        RECT 66.655 55.640 66.975 55.960 ;
        RECT 67.055 55.640 67.375 55.960 ;
        RECT 88.050 55.640 88.370 55.960 ;
        RECT 88.450 55.640 88.770 55.960 ;
        RECT 88.850 55.640 89.170 55.960 ;
        RECT 89.250 55.640 89.570 55.960 ;
        RECT 110.245 55.640 110.565 55.960 ;
        RECT 110.645 55.640 110.965 55.960 ;
        RECT 111.045 55.640 111.365 55.960 ;
        RECT 111.445 55.640 111.765 55.960 ;
        RECT 132.440 55.640 132.760 55.960 ;
        RECT 132.840 55.640 133.160 55.960 ;
        RECT 133.240 55.640 133.560 55.960 ;
        RECT 133.640 55.640 133.960 55.960 ;
        RECT 65.855 50.200 66.175 50.520 ;
        RECT 66.255 50.200 66.575 50.520 ;
        RECT 66.655 50.200 66.975 50.520 ;
        RECT 67.055 50.200 67.375 50.520 ;
        RECT 88.050 50.200 88.370 50.520 ;
        RECT 88.450 50.200 88.770 50.520 ;
        RECT 88.850 50.200 89.170 50.520 ;
        RECT 89.250 50.200 89.570 50.520 ;
        RECT 110.245 50.200 110.565 50.520 ;
        RECT 110.645 50.200 110.965 50.520 ;
        RECT 111.045 50.200 111.365 50.520 ;
        RECT 111.445 50.200 111.765 50.520 ;
        RECT 132.440 50.200 132.760 50.520 ;
        RECT 132.840 50.200 133.160 50.520 ;
        RECT 133.240 50.200 133.560 50.520 ;
        RECT 133.640 50.200 133.960 50.520 ;
        RECT 65.855 44.760 66.175 45.080 ;
        RECT 66.255 44.760 66.575 45.080 ;
        RECT 66.655 44.760 66.975 45.080 ;
        RECT 67.055 44.760 67.375 45.080 ;
        RECT 88.050 44.760 88.370 45.080 ;
        RECT 88.450 44.760 88.770 45.080 ;
        RECT 88.850 44.760 89.170 45.080 ;
        RECT 89.250 44.760 89.570 45.080 ;
        RECT 110.245 44.760 110.565 45.080 ;
        RECT 110.645 44.760 110.965 45.080 ;
        RECT 111.045 44.760 111.365 45.080 ;
        RECT 111.445 44.760 111.765 45.080 ;
        RECT 132.440 44.760 132.760 45.080 ;
        RECT 132.840 44.760 133.160 45.080 ;
        RECT 133.240 44.760 133.560 45.080 ;
        RECT 133.640 44.760 133.960 45.080 ;
        RECT 65.855 39.320 66.175 39.640 ;
        RECT 66.255 39.320 66.575 39.640 ;
        RECT 66.655 39.320 66.975 39.640 ;
        RECT 67.055 39.320 67.375 39.640 ;
        RECT 88.050 39.320 88.370 39.640 ;
        RECT 88.450 39.320 88.770 39.640 ;
        RECT 88.850 39.320 89.170 39.640 ;
        RECT 89.250 39.320 89.570 39.640 ;
        RECT 110.245 39.320 110.565 39.640 ;
        RECT 110.645 39.320 110.965 39.640 ;
        RECT 111.045 39.320 111.365 39.640 ;
        RECT 111.445 39.320 111.765 39.640 ;
        RECT 132.440 39.320 132.760 39.640 ;
        RECT 132.840 39.320 133.160 39.640 ;
        RECT 133.240 39.320 133.560 39.640 ;
        RECT 133.640 39.320 133.960 39.640 ;
        RECT 65.855 33.880 66.175 34.200 ;
        RECT 66.255 33.880 66.575 34.200 ;
        RECT 66.655 33.880 66.975 34.200 ;
        RECT 67.055 33.880 67.375 34.200 ;
        RECT 88.050 33.880 88.370 34.200 ;
        RECT 88.450 33.880 88.770 34.200 ;
        RECT 88.850 33.880 89.170 34.200 ;
        RECT 89.250 33.880 89.570 34.200 ;
        RECT 110.245 33.880 110.565 34.200 ;
        RECT 110.645 33.880 110.965 34.200 ;
        RECT 111.045 33.880 111.365 34.200 ;
        RECT 111.445 33.880 111.765 34.200 ;
        RECT 132.440 33.880 132.760 34.200 ;
        RECT 132.840 33.880 133.160 34.200 ;
        RECT 133.240 33.880 133.560 34.200 ;
        RECT 133.640 33.880 133.960 34.200 ;
        RECT 65.855 28.440 66.175 28.760 ;
        RECT 66.255 28.440 66.575 28.760 ;
        RECT 66.655 28.440 66.975 28.760 ;
        RECT 67.055 28.440 67.375 28.760 ;
        RECT 88.050 28.440 88.370 28.760 ;
        RECT 88.450 28.440 88.770 28.760 ;
        RECT 88.850 28.440 89.170 28.760 ;
        RECT 89.250 28.440 89.570 28.760 ;
        RECT 110.245 28.440 110.565 28.760 ;
        RECT 110.645 28.440 110.965 28.760 ;
        RECT 111.045 28.440 111.365 28.760 ;
        RECT 111.445 28.440 111.765 28.760 ;
        RECT 132.440 28.440 132.760 28.760 ;
        RECT 132.840 28.440 133.160 28.760 ;
        RECT 133.240 28.440 133.560 28.760 ;
        RECT 133.640 28.440 133.960 28.760 ;
      LAYER met4 ;
        RECT 65.815 25.640 67.415 102.280 ;
        RECT 88.010 25.640 89.610 102.280 ;
        RECT 110.205 25.640 111.805 102.280 ;
        RECT 132.400 25.640 134.000 102.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 68.545 101.195 68.715 101.720 ;
        RECT 81.425 101.195 81.595 101.720 ;
        RECT 94.305 101.195 94.475 101.720 ;
        RECT 107.185 101.195 107.355 101.720 ;
        RECT 120.065 101.195 120.235 101.720 ;
        RECT 132.945 101.195 133.115 101.720 ;
        RECT 68.545 96.920 68.715 97.445 ;
        RECT 94.305 96.920 94.475 97.445 ;
        RECT 120.065 96.920 120.235 97.445 ;
        RECT 81.425 95.755 81.595 96.280 ;
        RECT 107.185 95.755 107.355 96.280 ;
        RECT 132.945 95.755 133.115 96.280 ;
        RECT 68.545 91.480 68.715 92.005 ;
        RECT 94.305 91.480 94.475 92.005 ;
        RECT 120.065 91.480 120.235 92.005 ;
        RECT 81.425 90.315 81.595 90.840 ;
        RECT 107.185 90.315 107.355 90.840 ;
        RECT 132.945 90.315 133.115 90.840 ;
        RECT 68.545 86.040 68.715 86.565 ;
        RECT 94.305 86.040 94.475 86.565 ;
        RECT 120.065 86.040 120.235 86.565 ;
        RECT 81.425 84.875 81.595 85.400 ;
        RECT 107.185 84.875 107.355 85.400 ;
        RECT 132.945 84.875 133.115 85.400 ;
        RECT 68.545 80.600 68.715 81.125 ;
        RECT 94.305 80.600 94.475 81.125 ;
        RECT 120.065 80.600 120.235 81.125 ;
        RECT 81.425 79.435 81.595 79.960 ;
        RECT 107.185 79.435 107.355 79.960 ;
        RECT 132.945 79.435 133.115 79.960 ;
        RECT 68.545 75.160 68.715 75.685 ;
        RECT 94.305 75.160 94.475 75.685 ;
        RECT 120.065 75.160 120.235 75.685 ;
        RECT 81.425 73.995 81.595 74.520 ;
        RECT 107.185 73.995 107.355 74.520 ;
        RECT 132.945 73.995 133.115 74.520 ;
        RECT 68.545 69.720 68.715 70.245 ;
        RECT 94.305 69.720 94.475 70.245 ;
        RECT 120.065 69.720 120.235 70.245 ;
        RECT 81.425 68.555 81.595 69.080 ;
        RECT 107.185 68.555 107.355 69.080 ;
        RECT 132.945 68.555 133.115 69.080 ;
        RECT 68.545 64.280 68.715 64.805 ;
        RECT 94.305 64.280 94.475 64.805 ;
        RECT 120.065 64.280 120.235 64.805 ;
        RECT 81.425 63.115 81.595 63.640 ;
        RECT 107.185 63.115 107.355 63.640 ;
        RECT 132.945 63.115 133.115 63.640 ;
        RECT 68.545 58.840 68.715 59.365 ;
        RECT 94.305 58.840 94.475 59.365 ;
        RECT 120.065 58.840 120.235 59.365 ;
        RECT 81.425 57.675 81.595 58.200 ;
        RECT 107.185 57.675 107.355 58.200 ;
        RECT 132.945 57.675 133.115 58.200 ;
        RECT 68.545 53.400 68.715 53.925 ;
        RECT 94.305 53.400 94.475 53.925 ;
        RECT 120.065 53.400 120.235 53.925 ;
        RECT 81.425 52.235 81.595 52.760 ;
        RECT 107.185 52.235 107.355 52.760 ;
        RECT 132.945 52.235 133.115 52.760 ;
        RECT 68.545 47.960 68.715 48.485 ;
        RECT 94.305 47.960 94.475 48.485 ;
        RECT 120.065 47.960 120.235 48.485 ;
        RECT 81.425 46.795 81.595 47.320 ;
        RECT 107.185 46.795 107.355 47.320 ;
        RECT 132.945 46.795 133.115 47.320 ;
        RECT 68.545 42.520 68.715 43.045 ;
        RECT 94.305 42.520 94.475 43.045 ;
        RECT 120.065 42.520 120.235 43.045 ;
        RECT 81.425 41.355 81.595 41.880 ;
        RECT 107.185 41.355 107.355 41.880 ;
        RECT 132.945 41.355 133.115 41.880 ;
        RECT 68.545 37.080 68.715 37.605 ;
        RECT 94.305 37.080 94.475 37.605 ;
        RECT 120.065 37.080 120.235 37.605 ;
        RECT 81.425 35.915 81.595 36.440 ;
        RECT 107.185 35.915 107.355 36.440 ;
        RECT 132.945 35.915 133.115 36.440 ;
        RECT 68.545 31.640 68.715 32.165 ;
        RECT 94.305 31.640 94.475 32.165 ;
        RECT 120.065 31.640 120.235 32.165 ;
        RECT 81.425 30.475 81.595 31.000 ;
        RECT 107.185 30.475 107.355 31.000 ;
        RECT 132.945 30.475 133.115 31.000 ;
        RECT 68.545 26.200 68.715 26.725 ;
        RECT 81.425 26.200 81.595 26.725 ;
        RECT 94.305 26.200 94.475 26.725 ;
        RECT 107.185 26.200 107.355 26.725 ;
        RECT 120.065 26.200 120.235 26.725 ;
        RECT 132.945 26.200 133.115 26.725 ;
      LAYER li1 ;
        RECT 55.520 101.955 144.300 102.125 ;
        RECT 55.605 101.205 56.815 101.955 ;
        RECT 56.985 101.410 62.330 101.955 ;
        RECT 62.505 101.410 67.850 101.955 ;
        RECT 55.605 100.665 56.125 101.205 ;
        RECT 58.570 100.580 58.910 101.410 ;
        RECT 64.090 100.580 64.430 101.410 ;
        RECT 68.485 101.230 68.775 101.955 ;
        RECT 68.945 101.410 74.290 101.955 ;
        RECT 74.465 101.410 79.810 101.955 ;
        RECT 70.530 100.580 70.870 101.410 ;
        RECT 76.050 100.580 76.390 101.410 ;
        RECT 79.985 101.205 81.195 101.955 ;
        RECT 81.365 101.230 81.655 101.955 ;
        RECT 81.825 101.410 87.170 101.955 ;
        RECT 87.345 101.410 92.690 101.955 ;
        RECT 79.985 100.665 80.505 101.205 ;
        RECT 83.410 100.580 83.750 101.410 ;
        RECT 88.930 100.580 89.270 101.410 ;
        RECT 92.865 101.205 94.075 101.955 ;
        RECT 94.245 101.230 94.535 101.955 ;
        RECT 94.705 101.410 100.050 101.955 ;
        RECT 100.225 101.410 105.570 101.955 ;
        RECT 92.865 100.665 93.385 101.205 ;
        RECT 96.290 100.580 96.630 101.410 ;
        RECT 101.810 100.580 102.150 101.410 ;
        RECT 105.745 101.205 106.955 101.955 ;
        RECT 107.125 101.230 107.415 101.955 ;
        RECT 107.585 101.410 112.930 101.955 ;
        RECT 113.105 101.410 118.450 101.955 ;
        RECT 105.745 100.665 106.265 101.205 ;
        RECT 109.170 100.580 109.510 101.410 ;
        RECT 114.690 100.580 115.030 101.410 ;
        RECT 118.625 101.205 119.835 101.955 ;
        RECT 120.005 101.230 120.295 101.955 ;
        RECT 120.465 101.410 125.810 101.955 ;
        RECT 125.985 101.410 131.330 101.955 ;
        RECT 118.625 100.665 119.145 101.205 ;
        RECT 122.050 100.580 122.390 101.410 ;
        RECT 127.570 100.580 127.910 101.410 ;
        RECT 131.505 101.205 132.715 101.955 ;
        RECT 132.885 101.230 133.175 101.955 ;
        RECT 133.345 101.410 138.690 101.955 ;
        RECT 131.505 100.665 132.025 101.205 ;
        RECT 134.930 100.580 135.270 101.410 ;
        RECT 138.865 101.185 142.375 101.955 ;
        RECT 143.005 101.205 144.215 101.955 ;
        RECT 138.865 100.665 140.515 101.185 ;
        RECT 143.695 100.665 144.215 101.205 ;
        RECT 55.605 97.435 56.125 97.975 ;
        RECT 55.605 96.685 56.815 97.435 ;
        RECT 58.570 97.230 58.910 98.060 ;
        RECT 64.090 97.230 64.430 98.060 ;
        RECT 56.985 96.685 62.330 97.230 ;
        RECT 62.505 96.685 67.850 97.230 ;
        RECT 68.485 96.685 68.775 97.410 ;
        RECT 70.530 97.230 70.870 98.060 ;
        RECT 76.050 97.230 76.390 98.060 ;
        RECT 81.570 97.230 81.910 98.060 ;
        RECT 87.090 97.230 87.430 98.060 ;
        RECT 91.025 97.455 92.235 97.975 ;
        RECT 68.945 96.685 74.290 97.230 ;
        RECT 74.465 96.685 79.810 97.230 ;
        RECT 79.985 96.685 85.330 97.230 ;
        RECT 85.505 96.685 90.850 97.230 ;
        RECT 91.025 96.685 93.615 97.455 ;
        RECT 94.245 96.685 94.535 97.410 ;
        RECT 96.290 97.230 96.630 98.060 ;
        RECT 101.810 97.230 102.150 98.060 ;
        RECT 107.330 97.230 107.670 98.060 ;
        RECT 112.850 97.230 113.190 98.060 ;
        RECT 116.785 97.455 117.995 97.975 ;
        RECT 94.705 96.685 100.050 97.230 ;
        RECT 100.225 96.685 105.570 97.230 ;
        RECT 105.745 96.685 111.090 97.230 ;
        RECT 111.265 96.685 116.610 97.230 ;
        RECT 116.785 96.685 119.375 97.455 ;
        RECT 120.005 96.685 120.295 97.410 ;
        RECT 122.050 97.230 122.390 98.060 ;
        RECT 127.570 97.230 127.910 98.060 ;
        RECT 133.090 97.230 133.430 98.060 ;
        RECT 138.610 97.230 138.950 98.060 ;
        RECT 143.695 97.435 144.215 97.975 ;
        RECT 120.465 96.685 125.810 97.230 ;
        RECT 125.985 96.685 131.330 97.230 ;
        RECT 131.505 96.685 136.850 97.230 ;
        RECT 137.025 96.685 142.370 97.230 ;
        RECT 143.005 96.685 144.215 97.435 ;
        RECT 55.520 96.515 144.300 96.685 ;
        RECT 55.605 95.765 56.815 96.515 ;
        RECT 56.985 95.970 62.330 96.515 ;
        RECT 62.505 95.970 67.850 96.515 ;
        RECT 68.025 95.970 73.370 96.515 ;
        RECT 73.545 95.970 78.890 96.515 ;
        RECT 55.605 95.225 56.125 95.765 ;
        RECT 58.570 95.140 58.910 95.970 ;
        RECT 64.090 95.140 64.430 95.970 ;
        RECT 69.610 95.140 69.950 95.970 ;
        RECT 75.130 95.140 75.470 95.970 ;
        RECT 79.065 95.745 80.735 96.515 ;
        RECT 81.365 95.790 81.655 96.515 ;
        RECT 81.825 95.970 87.170 96.515 ;
        RECT 87.345 95.970 92.690 96.515 ;
        RECT 92.865 95.970 98.210 96.515 ;
        RECT 98.385 95.970 103.730 96.515 ;
        RECT 79.065 95.225 79.815 95.745 ;
        RECT 83.410 95.140 83.750 95.970 ;
        RECT 88.930 95.140 89.270 95.970 ;
        RECT 94.450 95.140 94.790 95.970 ;
        RECT 99.970 95.140 100.310 95.970 ;
        RECT 103.905 95.745 106.495 96.515 ;
        RECT 107.125 95.790 107.415 96.515 ;
        RECT 107.585 95.970 112.930 96.515 ;
        RECT 113.105 95.970 118.450 96.515 ;
        RECT 118.625 95.970 123.970 96.515 ;
        RECT 124.145 95.970 129.490 96.515 ;
        RECT 103.905 95.225 105.115 95.745 ;
        RECT 109.170 95.140 109.510 95.970 ;
        RECT 114.690 95.140 115.030 95.970 ;
        RECT 120.210 95.140 120.550 95.970 ;
        RECT 125.730 95.140 126.070 95.970 ;
        RECT 129.665 95.745 132.255 96.515 ;
        RECT 132.885 95.790 133.175 96.515 ;
        RECT 133.345 95.970 138.690 96.515 ;
        RECT 129.665 95.225 130.875 95.745 ;
        RECT 134.930 95.140 135.270 95.970 ;
        RECT 138.865 95.745 142.375 96.515 ;
        RECT 143.005 95.765 144.215 96.515 ;
        RECT 138.865 95.225 140.515 95.745 ;
        RECT 143.695 95.225 144.215 95.765 ;
        RECT 55.605 91.995 56.125 92.535 ;
        RECT 55.605 91.245 56.815 91.995 ;
        RECT 58.570 91.790 58.910 92.620 ;
        RECT 64.090 91.790 64.430 92.620 ;
        RECT 56.985 91.245 62.330 91.790 ;
        RECT 62.505 91.245 67.850 91.790 ;
        RECT 68.485 91.245 68.775 91.970 ;
        RECT 70.530 91.790 70.870 92.620 ;
        RECT 76.050 91.790 76.390 92.620 ;
        RECT 81.570 91.790 81.910 92.620 ;
        RECT 87.090 91.790 87.430 92.620 ;
        RECT 91.025 92.015 92.235 92.535 ;
        RECT 68.945 91.245 74.290 91.790 ;
        RECT 74.465 91.245 79.810 91.790 ;
        RECT 79.985 91.245 85.330 91.790 ;
        RECT 85.505 91.245 90.850 91.790 ;
        RECT 91.025 91.245 93.615 92.015 ;
        RECT 94.245 91.245 94.535 91.970 ;
        RECT 96.290 91.790 96.630 92.620 ;
        RECT 101.810 91.790 102.150 92.620 ;
        RECT 107.330 91.790 107.670 92.620 ;
        RECT 112.850 91.790 113.190 92.620 ;
        RECT 116.785 92.015 117.995 92.535 ;
        RECT 94.705 91.245 100.050 91.790 ;
        RECT 100.225 91.245 105.570 91.790 ;
        RECT 105.745 91.245 111.090 91.790 ;
        RECT 111.265 91.245 116.610 91.790 ;
        RECT 116.785 91.245 119.375 92.015 ;
        RECT 120.005 91.245 120.295 91.970 ;
        RECT 122.050 91.790 122.390 92.620 ;
        RECT 127.570 91.790 127.910 92.620 ;
        RECT 133.090 91.790 133.430 92.620 ;
        RECT 138.610 91.790 138.950 92.620 ;
        RECT 143.695 91.995 144.215 92.535 ;
        RECT 120.465 91.245 125.810 91.790 ;
        RECT 125.985 91.245 131.330 91.790 ;
        RECT 131.505 91.245 136.850 91.790 ;
        RECT 137.025 91.245 142.370 91.790 ;
        RECT 143.005 91.245 144.215 91.995 ;
        RECT 55.520 91.075 144.300 91.245 ;
        RECT 55.605 90.325 56.815 91.075 ;
        RECT 56.985 90.530 62.330 91.075 ;
        RECT 62.505 90.530 67.850 91.075 ;
        RECT 68.025 90.530 73.370 91.075 ;
        RECT 73.545 90.530 78.890 91.075 ;
        RECT 55.605 89.785 56.125 90.325 ;
        RECT 58.570 89.700 58.910 90.530 ;
        RECT 64.090 89.700 64.430 90.530 ;
        RECT 69.610 89.700 69.950 90.530 ;
        RECT 75.130 89.700 75.470 90.530 ;
        RECT 79.065 90.305 80.735 91.075 ;
        RECT 81.365 90.350 81.655 91.075 ;
        RECT 81.825 90.530 87.170 91.075 ;
        RECT 87.345 90.530 92.690 91.075 ;
        RECT 92.865 90.530 98.210 91.075 ;
        RECT 98.385 90.530 103.730 91.075 ;
        RECT 79.065 89.785 79.815 90.305 ;
        RECT 83.410 89.700 83.750 90.530 ;
        RECT 88.930 89.700 89.270 90.530 ;
        RECT 94.450 89.700 94.790 90.530 ;
        RECT 99.970 89.700 100.310 90.530 ;
        RECT 103.905 90.305 106.495 91.075 ;
        RECT 107.125 90.350 107.415 91.075 ;
        RECT 107.585 90.530 112.930 91.075 ;
        RECT 113.105 90.530 118.450 91.075 ;
        RECT 118.625 90.530 123.970 91.075 ;
        RECT 124.145 90.530 129.490 91.075 ;
        RECT 103.905 89.785 105.115 90.305 ;
        RECT 109.170 89.700 109.510 90.530 ;
        RECT 114.690 89.700 115.030 90.530 ;
        RECT 120.210 89.700 120.550 90.530 ;
        RECT 125.730 89.700 126.070 90.530 ;
        RECT 129.665 90.305 132.255 91.075 ;
        RECT 132.885 90.350 133.175 91.075 ;
        RECT 133.345 90.530 138.690 91.075 ;
        RECT 129.665 89.785 130.875 90.305 ;
        RECT 134.930 89.700 135.270 90.530 ;
        RECT 138.865 90.305 142.375 91.075 ;
        RECT 143.005 90.325 144.215 91.075 ;
        RECT 138.865 89.785 140.515 90.305 ;
        RECT 143.695 89.785 144.215 90.325 ;
        RECT 55.605 86.555 56.125 87.095 ;
        RECT 55.605 85.805 56.815 86.555 ;
        RECT 58.570 86.350 58.910 87.180 ;
        RECT 64.090 86.350 64.430 87.180 ;
        RECT 56.985 85.805 62.330 86.350 ;
        RECT 62.505 85.805 67.850 86.350 ;
        RECT 68.485 85.805 68.775 86.530 ;
        RECT 70.530 86.350 70.870 87.180 ;
        RECT 76.050 86.350 76.390 87.180 ;
        RECT 81.570 86.350 81.910 87.180 ;
        RECT 87.090 86.350 87.430 87.180 ;
        RECT 91.025 86.575 92.235 87.095 ;
        RECT 68.945 85.805 74.290 86.350 ;
        RECT 74.465 85.805 79.810 86.350 ;
        RECT 79.985 85.805 85.330 86.350 ;
        RECT 85.505 85.805 90.850 86.350 ;
        RECT 91.025 85.805 93.615 86.575 ;
        RECT 94.245 85.805 94.535 86.530 ;
        RECT 96.290 86.350 96.630 87.180 ;
        RECT 101.810 86.350 102.150 87.180 ;
        RECT 107.330 86.350 107.670 87.180 ;
        RECT 112.850 86.350 113.190 87.180 ;
        RECT 116.785 86.575 117.995 87.095 ;
        RECT 94.705 85.805 100.050 86.350 ;
        RECT 100.225 85.805 105.570 86.350 ;
        RECT 105.745 85.805 111.090 86.350 ;
        RECT 111.265 85.805 116.610 86.350 ;
        RECT 116.785 85.805 119.375 86.575 ;
        RECT 120.005 85.805 120.295 86.530 ;
        RECT 122.050 86.350 122.390 87.180 ;
        RECT 127.570 86.350 127.910 87.180 ;
        RECT 133.090 86.350 133.430 87.180 ;
        RECT 138.610 86.350 138.950 87.180 ;
        RECT 143.695 86.555 144.215 87.095 ;
        RECT 120.465 85.805 125.810 86.350 ;
        RECT 125.985 85.805 131.330 86.350 ;
        RECT 131.505 85.805 136.850 86.350 ;
        RECT 137.025 85.805 142.370 86.350 ;
        RECT 143.005 85.805 144.215 86.555 ;
        RECT 55.520 85.635 144.300 85.805 ;
        RECT 55.605 84.885 56.815 85.635 ;
        RECT 56.985 85.090 62.330 85.635 ;
        RECT 62.505 85.090 67.850 85.635 ;
        RECT 68.025 85.090 73.370 85.635 ;
        RECT 73.545 85.090 78.890 85.635 ;
        RECT 55.605 84.345 56.125 84.885 ;
        RECT 58.570 84.260 58.910 85.090 ;
        RECT 64.090 84.260 64.430 85.090 ;
        RECT 69.610 84.260 69.950 85.090 ;
        RECT 75.130 84.260 75.470 85.090 ;
        RECT 79.065 84.865 80.735 85.635 ;
        RECT 81.365 84.910 81.655 85.635 ;
        RECT 81.825 85.090 87.170 85.635 ;
        RECT 87.345 85.090 92.690 85.635 ;
        RECT 92.865 85.090 98.210 85.635 ;
        RECT 98.385 85.090 103.730 85.635 ;
        RECT 79.065 84.345 79.815 84.865 ;
        RECT 83.410 84.260 83.750 85.090 ;
        RECT 88.930 84.260 89.270 85.090 ;
        RECT 94.450 84.260 94.790 85.090 ;
        RECT 99.970 84.260 100.310 85.090 ;
        RECT 103.905 84.865 106.495 85.635 ;
        RECT 107.125 84.910 107.415 85.635 ;
        RECT 107.585 85.090 112.930 85.635 ;
        RECT 113.105 85.090 118.450 85.635 ;
        RECT 118.625 85.090 123.970 85.635 ;
        RECT 124.145 85.090 129.490 85.635 ;
        RECT 103.905 84.345 105.115 84.865 ;
        RECT 109.170 84.260 109.510 85.090 ;
        RECT 114.690 84.260 115.030 85.090 ;
        RECT 120.210 84.260 120.550 85.090 ;
        RECT 125.730 84.260 126.070 85.090 ;
        RECT 129.665 84.865 132.255 85.635 ;
        RECT 132.885 84.910 133.175 85.635 ;
        RECT 133.345 85.090 138.690 85.635 ;
        RECT 129.665 84.345 130.875 84.865 ;
        RECT 134.930 84.260 135.270 85.090 ;
        RECT 138.865 84.865 142.375 85.635 ;
        RECT 143.005 84.885 144.215 85.635 ;
        RECT 138.865 84.345 140.515 84.865 ;
        RECT 143.695 84.345 144.215 84.885 ;
        RECT 55.605 81.115 56.125 81.655 ;
        RECT 55.605 80.365 56.815 81.115 ;
        RECT 58.570 80.910 58.910 81.740 ;
        RECT 64.090 80.910 64.430 81.740 ;
        RECT 56.985 80.365 62.330 80.910 ;
        RECT 62.505 80.365 67.850 80.910 ;
        RECT 68.485 80.365 68.775 81.090 ;
        RECT 70.530 80.910 70.870 81.740 ;
        RECT 76.050 80.910 76.390 81.740 ;
        RECT 81.570 80.910 81.910 81.740 ;
        RECT 87.090 80.910 87.430 81.740 ;
        RECT 91.025 81.135 92.235 81.655 ;
        RECT 68.945 80.365 74.290 80.910 ;
        RECT 74.465 80.365 79.810 80.910 ;
        RECT 79.985 80.365 85.330 80.910 ;
        RECT 85.505 80.365 90.850 80.910 ;
        RECT 91.025 80.365 93.615 81.135 ;
        RECT 94.245 80.365 94.535 81.090 ;
        RECT 96.290 80.910 96.630 81.740 ;
        RECT 101.810 80.910 102.150 81.740 ;
        RECT 107.330 80.910 107.670 81.740 ;
        RECT 112.850 80.910 113.190 81.740 ;
        RECT 116.785 81.135 117.995 81.655 ;
        RECT 94.705 80.365 100.050 80.910 ;
        RECT 100.225 80.365 105.570 80.910 ;
        RECT 105.745 80.365 111.090 80.910 ;
        RECT 111.265 80.365 116.610 80.910 ;
        RECT 116.785 80.365 119.375 81.135 ;
        RECT 120.005 80.365 120.295 81.090 ;
        RECT 122.050 80.910 122.390 81.740 ;
        RECT 127.570 80.910 127.910 81.740 ;
        RECT 133.090 80.910 133.430 81.740 ;
        RECT 138.610 80.910 138.950 81.740 ;
        RECT 143.695 81.115 144.215 81.655 ;
        RECT 120.465 80.365 125.810 80.910 ;
        RECT 125.985 80.365 131.330 80.910 ;
        RECT 131.505 80.365 136.850 80.910 ;
        RECT 137.025 80.365 142.370 80.910 ;
        RECT 143.005 80.365 144.215 81.115 ;
        RECT 55.520 80.195 144.300 80.365 ;
        RECT 55.605 79.445 56.815 80.195 ;
        RECT 56.985 79.650 62.330 80.195 ;
        RECT 62.505 79.650 67.850 80.195 ;
        RECT 68.025 79.650 73.370 80.195 ;
        RECT 73.545 79.650 78.890 80.195 ;
        RECT 55.605 78.905 56.125 79.445 ;
        RECT 58.570 78.820 58.910 79.650 ;
        RECT 64.090 78.820 64.430 79.650 ;
        RECT 69.610 78.820 69.950 79.650 ;
        RECT 75.130 78.820 75.470 79.650 ;
        RECT 79.065 79.425 80.735 80.195 ;
        RECT 81.365 79.470 81.655 80.195 ;
        RECT 81.825 79.650 87.170 80.195 ;
        RECT 87.345 79.650 92.690 80.195 ;
        RECT 92.865 79.650 98.210 80.195 ;
        RECT 98.385 79.650 103.730 80.195 ;
        RECT 79.065 78.905 79.815 79.425 ;
        RECT 83.410 78.820 83.750 79.650 ;
        RECT 88.930 78.820 89.270 79.650 ;
        RECT 94.450 78.820 94.790 79.650 ;
        RECT 99.970 78.820 100.310 79.650 ;
        RECT 103.905 79.425 106.495 80.195 ;
        RECT 107.125 79.470 107.415 80.195 ;
        RECT 107.585 79.650 112.930 80.195 ;
        RECT 113.105 79.650 118.450 80.195 ;
        RECT 118.625 79.650 123.970 80.195 ;
        RECT 124.145 79.650 129.490 80.195 ;
        RECT 103.905 78.905 105.115 79.425 ;
        RECT 109.170 78.820 109.510 79.650 ;
        RECT 114.690 78.820 115.030 79.650 ;
        RECT 120.210 78.820 120.550 79.650 ;
        RECT 125.730 78.820 126.070 79.650 ;
        RECT 129.665 79.425 132.255 80.195 ;
        RECT 132.885 79.470 133.175 80.195 ;
        RECT 133.345 79.650 138.690 80.195 ;
        RECT 129.665 78.905 130.875 79.425 ;
        RECT 134.930 78.820 135.270 79.650 ;
        RECT 138.865 79.425 142.375 80.195 ;
        RECT 143.005 79.445 144.215 80.195 ;
        RECT 138.865 78.905 140.515 79.425 ;
        RECT 143.695 78.905 144.215 79.445 ;
        RECT 55.605 75.675 56.125 76.215 ;
        RECT 55.605 74.925 56.815 75.675 ;
        RECT 58.570 75.470 58.910 76.300 ;
        RECT 64.090 75.470 64.430 76.300 ;
        RECT 56.985 74.925 62.330 75.470 ;
        RECT 62.505 74.925 67.850 75.470 ;
        RECT 68.485 74.925 68.775 75.650 ;
        RECT 70.530 75.470 70.870 76.300 ;
        RECT 76.050 75.470 76.390 76.300 ;
        RECT 81.570 75.470 81.910 76.300 ;
        RECT 87.090 75.470 87.430 76.300 ;
        RECT 91.025 75.695 92.235 76.215 ;
        RECT 68.945 74.925 74.290 75.470 ;
        RECT 74.465 74.925 79.810 75.470 ;
        RECT 79.985 74.925 85.330 75.470 ;
        RECT 85.505 74.925 90.850 75.470 ;
        RECT 91.025 74.925 93.615 75.695 ;
        RECT 94.245 74.925 94.535 75.650 ;
        RECT 96.290 75.470 96.630 76.300 ;
        RECT 101.810 75.470 102.150 76.300 ;
        RECT 107.330 75.470 107.670 76.300 ;
        RECT 112.850 75.470 113.190 76.300 ;
        RECT 116.785 75.695 117.995 76.215 ;
        RECT 94.705 74.925 100.050 75.470 ;
        RECT 100.225 74.925 105.570 75.470 ;
        RECT 105.745 74.925 111.090 75.470 ;
        RECT 111.265 74.925 116.610 75.470 ;
        RECT 116.785 74.925 119.375 75.695 ;
        RECT 120.005 74.925 120.295 75.650 ;
        RECT 122.050 75.470 122.390 76.300 ;
        RECT 127.570 75.470 127.910 76.300 ;
        RECT 133.090 75.470 133.430 76.300 ;
        RECT 138.610 75.470 138.950 76.300 ;
        RECT 143.695 75.675 144.215 76.215 ;
        RECT 120.465 74.925 125.810 75.470 ;
        RECT 125.985 74.925 131.330 75.470 ;
        RECT 131.505 74.925 136.850 75.470 ;
        RECT 137.025 74.925 142.370 75.470 ;
        RECT 143.005 74.925 144.215 75.675 ;
        RECT 55.520 74.755 144.300 74.925 ;
        RECT 55.605 74.005 56.815 74.755 ;
        RECT 56.985 74.210 62.330 74.755 ;
        RECT 62.505 74.210 67.850 74.755 ;
        RECT 55.605 73.465 56.125 74.005 ;
        RECT 58.570 73.380 58.910 74.210 ;
        RECT 64.090 73.380 64.430 74.210 ;
        RECT 68.025 73.985 69.695 74.755 ;
        RECT 68.025 73.465 68.775 73.985 ;
        RECT 70.365 73.935 70.595 74.755 ;
        RECT 71.265 73.935 71.475 74.755 ;
        RECT 72.180 74.375 72.510 74.755 ;
        RECT 73.110 73.915 73.370 74.755 ;
        RECT 73.545 74.210 78.890 74.755 ;
        RECT 75.130 73.380 75.470 74.210 ;
        RECT 79.065 73.985 80.735 74.755 ;
        RECT 81.365 74.030 81.655 74.755 ;
        RECT 81.825 74.210 87.170 74.755 ;
        RECT 87.345 74.210 92.690 74.755 ;
        RECT 92.865 74.210 98.210 74.755 ;
        RECT 98.385 74.210 103.730 74.755 ;
        RECT 79.065 73.465 79.815 73.985 ;
        RECT 83.410 73.380 83.750 74.210 ;
        RECT 88.930 73.380 89.270 74.210 ;
        RECT 94.450 73.380 94.790 74.210 ;
        RECT 99.970 73.380 100.310 74.210 ;
        RECT 103.905 73.985 106.495 74.755 ;
        RECT 107.125 74.030 107.415 74.755 ;
        RECT 107.585 74.210 112.930 74.755 ;
        RECT 113.105 74.210 118.450 74.755 ;
        RECT 118.625 74.210 123.970 74.755 ;
        RECT 124.145 74.210 129.490 74.755 ;
        RECT 103.905 73.465 105.115 73.985 ;
        RECT 109.170 73.380 109.510 74.210 ;
        RECT 114.690 73.380 115.030 74.210 ;
        RECT 120.210 73.380 120.550 74.210 ;
        RECT 125.730 73.380 126.070 74.210 ;
        RECT 129.665 73.985 132.255 74.755 ;
        RECT 132.885 74.030 133.175 74.755 ;
        RECT 133.345 74.210 138.690 74.755 ;
        RECT 129.665 73.465 130.875 73.985 ;
        RECT 134.930 73.380 135.270 74.210 ;
        RECT 138.865 73.985 142.375 74.755 ;
        RECT 143.005 74.005 144.215 74.755 ;
        RECT 138.865 73.465 140.515 73.985 ;
        RECT 143.695 73.465 144.215 74.005 ;
        RECT 55.605 70.235 56.125 70.775 ;
        RECT 56.985 70.255 58.635 70.775 ;
        RECT 55.605 69.485 56.815 70.235 ;
        RECT 56.985 69.485 60.495 70.255 ;
        RECT 61.185 69.485 61.395 70.305 ;
        RECT 62.065 69.485 62.295 70.305 ;
        RECT 62.505 69.485 62.815 70.285 ;
        RECT 64.525 69.485 65.285 69.965 ;
        RECT 66.635 69.485 66.965 69.845 ;
        RECT 68.485 69.485 68.775 70.210 ;
        RECT 70.530 70.030 70.870 70.860 ;
        RECT 76.050 70.030 76.390 70.860 ;
        RECT 81.570 70.030 81.910 70.860 ;
        RECT 87.090 70.030 87.430 70.860 ;
        RECT 91.025 70.255 92.235 70.775 ;
        RECT 68.945 69.485 74.290 70.030 ;
        RECT 74.465 69.485 79.810 70.030 ;
        RECT 79.985 69.485 85.330 70.030 ;
        RECT 85.505 69.485 90.850 70.030 ;
        RECT 91.025 69.485 93.615 70.255 ;
        RECT 94.245 69.485 94.535 70.210 ;
        RECT 96.290 70.030 96.630 70.860 ;
        RECT 101.810 70.030 102.150 70.860 ;
        RECT 107.330 70.030 107.670 70.860 ;
        RECT 112.850 70.030 113.190 70.860 ;
        RECT 116.785 70.255 117.995 70.775 ;
        RECT 94.705 69.485 100.050 70.030 ;
        RECT 100.225 69.485 105.570 70.030 ;
        RECT 105.745 69.485 111.090 70.030 ;
        RECT 111.265 69.485 116.610 70.030 ;
        RECT 116.785 69.485 119.375 70.255 ;
        RECT 120.005 69.485 120.295 70.210 ;
        RECT 122.050 70.030 122.390 70.860 ;
        RECT 127.570 70.030 127.910 70.860 ;
        RECT 133.090 70.030 133.430 70.860 ;
        RECT 138.610 70.030 138.950 70.860 ;
        RECT 143.695 70.235 144.215 70.775 ;
        RECT 120.465 69.485 125.810 70.030 ;
        RECT 125.985 69.485 131.330 70.030 ;
        RECT 131.505 69.485 136.850 70.030 ;
        RECT 137.025 69.485 142.370 70.030 ;
        RECT 143.005 69.485 144.215 70.235 ;
        RECT 55.520 69.315 144.300 69.485 ;
        RECT 55.605 68.565 56.815 69.315 ;
        RECT 57.425 68.935 57.755 69.315 ;
        RECT 58.365 68.770 63.710 69.315 ;
        RECT 65.315 68.855 65.485 69.315 ;
        RECT 67.535 68.805 67.870 69.315 ;
        RECT 69.360 68.915 69.690 69.315 ;
        RECT 71.245 68.770 76.590 69.315 ;
        RECT 55.605 68.025 56.125 68.565 ;
        RECT 59.950 67.940 60.290 68.770 ;
        RECT 72.830 67.940 73.170 68.770 ;
        RECT 76.765 68.545 80.275 69.315 ;
        RECT 81.365 68.590 81.655 69.315 ;
        RECT 81.825 68.770 87.170 69.315 ;
        RECT 87.345 68.770 92.690 69.315 ;
        RECT 92.865 68.770 98.210 69.315 ;
        RECT 98.385 68.770 103.730 69.315 ;
        RECT 76.765 68.025 78.415 68.545 ;
        RECT 83.410 67.940 83.750 68.770 ;
        RECT 88.930 67.940 89.270 68.770 ;
        RECT 94.450 67.940 94.790 68.770 ;
        RECT 99.970 67.940 100.310 68.770 ;
        RECT 103.905 68.545 106.495 69.315 ;
        RECT 107.125 68.590 107.415 69.315 ;
        RECT 107.585 68.770 112.930 69.315 ;
        RECT 113.105 68.770 118.450 69.315 ;
        RECT 118.625 68.770 123.970 69.315 ;
        RECT 124.145 68.770 129.490 69.315 ;
        RECT 103.905 68.025 105.115 68.545 ;
        RECT 109.170 67.940 109.510 68.770 ;
        RECT 114.690 67.940 115.030 68.770 ;
        RECT 120.210 67.940 120.550 68.770 ;
        RECT 125.730 67.940 126.070 68.770 ;
        RECT 129.665 68.545 132.255 69.315 ;
        RECT 132.885 68.590 133.175 69.315 ;
        RECT 133.345 68.770 138.690 69.315 ;
        RECT 129.665 68.025 130.875 68.545 ;
        RECT 134.930 67.940 135.270 68.770 ;
        RECT 138.865 68.545 142.375 69.315 ;
        RECT 143.005 68.565 144.215 69.315 ;
        RECT 138.865 68.025 140.515 68.545 ;
        RECT 143.695 68.025 144.215 68.565 ;
        RECT 55.605 64.795 56.125 65.335 ;
        RECT 55.605 64.045 56.815 64.795 ;
        RECT 59.950 64.590 60.290 65.420 ;
        RECT 63.885 64.815 65.535 65.335 ;
        RECT 57.425 64.045 57.755 64.425 ;
        RECT 58.365 64.045 63.710 64.590 ;
        RECT 63.885 64.045 67.395 64.815 ;
        RECT 68.485 64.045 68.775 64.770 ;
        RECT 70.530 64.590 70.870 65.420 ;
        RECT 76.050 64.590 76.390 65.420 ;
        RECT 81.570 64.590 81.910 65.420 ;
        RECT 87.090 64.590 87.430 65.420 ;
        RECT 91.025 64.815 92.235 65.335 ;
        RECT 68.945 64.045 74.290 64.590 ;
        RECT 74.465 64.045 79.810 64.590 ;
        RECT 79.985 64.045 85.330 64.590 ;
        RECT 85.505 64.045 90.850 64.590 ;
        RECT 91.025 64.045 93.615 64.815 ;
        RECT 94.245 64.045 94.535 64.770 ;
        RECT 96.290 64.590 96.630 65.420 ;
        RECT 101.810 64.590 102.150 65.420 ;
        RECT 107.330 64.590 107.670 65.420 ;
        RECT 112.850 64.590 113.190 65.420 ;
        RECT 116.785 64.815 117.995 65.335 ;
        RECT 94.705 64.045 100.050 64.590 ;
        RECT 100.225 64.045 105.570 64.590 ;
        RECT 105.745 64.045 111.090 64.590 ;
        RECT 111.265 64.045 116.610 64.590 ;
        RECT 116.785 64.045 119.375 64.815 ;
        RECT 120.005 64.045 120.295 64.770 ;
        RECT 122.050 64.590 122.390 65.420 ;
        RECT 127.570 64.590 127.910 65.420 ;
        RECT 133.090 64.590 133.430 65.420 ;
        RECT 138.610 64.590 138.950 65.420 ;
        RECT 143.695 64.795 144.215 65.335 ;
        RECT 120.465 64.045 125.810 64.590 ;
        RECT 125.985 64.045 131.330 64.590 ;
        RECT 131.505 64.045 136.850 64.590 ;
        RECT 137.025 64.045 142.370 64.590 ;
        RECT 143.005 64.045 144.215 64.795 ;
        RECT 55.520 63.875 144.300 64.045 ;
        RECT 55.605 63.125 56.815 63.875 ;
        RECT 56.985 63.330 62.330 63.875 ;
        RECT 55.605 62.585 56.125 63.125 ;
        RECT 58.570 62.500 58.910 63.330 ;
        RECT 62.505 63.105 65.095 63.875 ;
        RECT 66.165 63.495 66.495 63.875 ;
        RECT 67.105 63.330 72.450 63.875 ;
        RECT 72.625 63.330 77.970 63.875 ;
        RECT 62.505 62.585 63.715 63.105 ;
        RECT 68.690 62.500 69.030 63.330 ;
        RECT 74.210 62.500 74.550 63.330 ;
        RECT 78.145 63.105 80.735 63.875 ;
        RECT 81.365 63.150 81.655 63.875 ;
        RECT 81.825 63.330 87.170 63.875 ;
        RECT 87.345 63.330 92.690 63.875 ;
        RECT 92.865 63.330 98.210 63.875 ;
        RECT 98.385 63.330 103.730 63.875 ;
        RECT 78.145 62.585 79.355 63.105 ;
        RECT 83.410 62.500 83.750 63.330 ;
        RECT 88.930 62.500 89.270 63.330 ;
        RECT 94.450 62.500 94.790 63.330 ;
        RECT 99.970 62.500 100.310 63.330 ;
        RECT 103.905 63.105 106.495 63.875 ;
        RECT 107.125 63.150 107.415 63.875 ;
        RECT 107.585 63.330 112.930 63.875 ;
        RECT 113.105 63.330 118.450 63.875 ;
        RECT 118.625 63.330 123.970 63.875 ;
        RECT 124.145 63.330 129.490 63.875 ;
        RECT 103.905 62.585 105.115 63.105 ;
        RECT 109.170 62.500 109.510 63.330 ;
        RECT 114.690 62.500 115.030 63.330 ;
        RECT 120.210 62.500 120.550 63.330 ;
        RECT 125.730 62.500 126.070 63.330 ;
        RECT 129.665 63.105 132.255 63.875 ;
        RECT 132.885 63.150 133.175 63.875 ;
        RECT 133.345 63.330 138.690 63.875 ;
        RECT 129.665 62.585 130.875 63.105 ;
        RECT 134.930 62.500 135.270 63.330 ;
        RECT 138.865 63.105 142.375 63.875 ;
        RECT 143.005 63.125 144.215 63.875 ;
        RECT 138.865 62.585 140.515 63.105 ;
        RECT 143.695 62.585 144.215 63.125 ;
        RECT 55.605 59.355 56.125 59.895 ;
        RECT 55.605 58.605 56.815 59.355 ;
        RECT 58.570 59.150 58.910 59.980 ;
        RECT 62.505 59.375 64.155 59.895 ;
        RECT 56.985 58.605 62.330 59.150 ;
        RECT 62.505 58.605 66.015 59.375 ;
        RECT 67.545 58.605 67.855 59.405 ;
        RECT 68.485 58.605 68.775 59.330 ;
        RECT 70.530 59.150 70.870 59.980 ;
        RECT 76.050 59.150 76.390 59.980 ;
        RECT 81.570 59.150 81.910 59.980 ;
        RECT 87.090 59.150 87.430 59.980 ;
        RECT 91.025 59.375 92.235 59.895 ;
        RECT 68.945 58.605 74.290 59.150 ;
        RECT 74.465 58.605 79.810 59.150 ;
        RECT 79.985 58.605 85.330 59.150 ;
        RECT 85.505 58.605 90.850 59.150 ;
        RECT 91.025 58.605 93.615 59.375 ;
        RECT 94.245 58.605 94.535 59.330 ;
        RECT 96.290 59.150 96.630 59.980 ;
        RECT 101.810 59.150 102.150 59.980 ;
        RECT 107.330 59.150 107.670 59.980 ;
        RECT 112.850 59.150 113.190 59.980 ;
        RECT 116.785 59.375 117.995 59.895 ;
        RECT 94.705 58.605 100.050 59.150 ;
        RECT 100.225 58.605 105.570 59.150 ;
        RECT 105.745 58.605 111.090 59.150 ;
        RECT 111.265 58.605 116.610 59.150 ;
        RECT 116.785 58.605 119.375 59.375 ;
        RECT 120.005 58.605 120.295 59.330 ;
        RECT 122.050 59.150 122.390 59.980 ;
        RECT 127.570 59.150 127.910 59.980 ;
        RECT 133.090 59.150 133.430 59.980 ;
        RECT 138.610 59.150 138.950 59.980 ;
        RECT 143.695 59.355 144.215 59.895 ;
        RECT 120.465 58.605 125.810 59.150 ;
        RECT 125.985 58.605 131.330 59.150 ;
        RECT 131.505 58.605 136.850 59.150 ;
        RECT 137.025 58.605 142.370 59.150 ;
        RECT 143.005 58.605 144.215 59.355 ;
        RECT 55.520 58.435 144.300 58.605 ;
        RECT 55.605 57.685 56.815 58.435 ;
        RECT 55.605 57.145 56.125 57.685 ;
        RECT 56.985 57.665 60.495 58.435 ;
        RECT 62.325 57.900 62.835 58.435 ;
        RECT 64.795 58.035 65.125 58.435 ;
        RECT 66.155 58.035 66.485 58.435 ;
        RECT 68.445 57.900 68.955 58.435 ;
        RECT 56.985 57.145 58.635 57.665 ;
        RECT 69.905 57.615 70.135 58.435 ;
        RECT 70.805 57.615 71.015 58.435 ;
        RECT 71.285 57.615 71.515 58.435 ;
        RECT 72.185 57.615 72.395 58.435 ;
        RECT 72.625 57.890 77.970 58.435 ;
        RECT 74.210 57.060 74.550 57.890 ;
        RECT 78.145 57.665 80.735 58.435 ;
        RECT 81.365 57.710 81.655 58.435 ;
        RECT 81.825 57.890 87.170 58.435 ;
        RECT 87.345 57.890 92.690 58.435 ;
        RECT 92.865 57.890 98.210 58.435 ;
        RECT 98.385 57.890 103.730 58.435 ;
        RECT 78.145 57.145 79.355 57.665 ;
        RECT 83.410 57.060 83.750 57.890 ;
        RECT 88.930 57.060 89.270 57.890 ;
        RECT 94.450 57.060 94.790 57.890 ;
        RECT 99.970 57.060 100.310 57.890 ;
        RECT 103.905 57.665 106.495 58.435 ;
        RECT 107.125 57.710 107.415 58.435 ;
        RECT 107.585 57.890 112.930 58.435 ;
        RECT 113.105 57.890 118.450 58.435 ;
        RECT 118.625 57.890 123.970 58.435 ;
        RECT 124.145 57.890 129.490 58.435 ;
        RECT 103.905 57.145 105.115 57.665 ;
        RECT 109.170 57.060 109.510 57.890 ;
        RECT 114.690 57.060 115.030 57.890 ;
        RECT 120.210 57.060 120.550 57.890 ;
        RECT 125.730 57.060 126.070 57.890 ;
        RECT 129.665 57.665 132.255 58.435 ;
        RECT 132.885 57.710 133.175 58.435 ;
        RECT 133.345 57.890 138.690 58.435 ;
        RECT 129.665 57.145 130.875 57.665 ;
        RECT 134.930 57.060 135.270 57.890 ;
        RECT 138.865 57.665 142.375 58.435 ;
        RECT 143.005 57.685 144.215 58.435 ;
        RECT 138.865 57.145 140.515 57.665 ;
        RECT 143.695 57.145 144.215 57.685 ;
        RECT 55.605 53.915 56.125 54.455 ;
        RECT 55.605 53.165 56.815 53.915 ;
        RECT 58.570 53.710 58.910 54.540 ;
        RECT 62.505 53.935 63.715 54.455 ;
        RECT 56.985 53.165 62.330 53.710 ;
        RECT 62.505 53.165 65.095 53.935 ;
        RECT 65.705 53.165 66.035 53.545 ;
        RECT 66.685 53.165 66.915 53.985 ;
        RECT 67.585 53.165 67.795 53.985 ;
        RECT 68.485 53.165 68.775 53.890 ;
        RECT 70.530 53.710 70.870 54.540 ;
        RECT 76.050 53.710 76.390 54.540 ;
        RECT 81.570 53.710 81.910 54.540 ;
        RECT 87.090 53.710 87.430 54.540 ;
        RECT 91.025 53.935 92.235 54.455 ;
        RECT 68.945 53.165 74.290 53.710 ;
        RECT 74.465 53.165 79.810 53.710 ;
        RECT 79.985 53.165 85.330 53.710 ;
        RECT 85.505 53.165 90.850 53.710 ;
        RECT 91.025 53.165 93.615 53.935 ;
        RECT 94.245 53.165 94.535 53.890 ;
        RECT 96.290 53.710 96.630 54.540 ;
        RECT 101.810 53.710 102.150 54.540 ;
        RECT 107.330 53.710 107.670 54.540 ;
        RECT 112.850 53.710 113.190 54.540 ;
        RECT 116.785 53.935 117.995 54.455 ;
        RECT 94.705 53.165 100.050 53.710 ;
        RECT 100.225 53.165 105.570 53.710 ;
        RECT 105.745 53.165 111.090 53.710 ;
        RECT 111.265 53.165 116.610 53.710 ;
        RECT 116.785 53.165 119.375 53.935 ;
        RECT 120.005 53.165 120.295 53.890 ;
        RECT 122.050 53.710 122.390 54.540 ;
        RECT 127.570 53.710 127.910 54.540 ;
        RECT 133.090 53.710 133.430 54.540 ;
        RECT 138.610 53.710 138.950 54.540 ;
        RECT 143.695 53.915 144.215 54.455 ;
        RECT 120.465 53.165 125.810 53.710 ;
        RECT 125.985 53.165 131.330 53.710 ;
        RECT 131.505 53.165 136.850 53.710 ;
        RECT 137.025 53.165 142.370 53.710 ;
        RECT 143.005 53.165 144.215 53.915 ;
        RECT 55.520 52.995 144.300 53.165 ;
        RECT 55.605 52.245 56.815 52.995 ;
        RECT 56.985 52.450 62.330 52.995 ;
        RECT 62.505 52.450 67.850 52.995 ;
        RECT 68.025 52.450 73.370 52.995 ;
        RECT 73.545 52.450 78.890 52.995 ;
        RECT 55.605 51.705 56.125 52.245 ;
        RECT 58.570 51.620 58.910 52.450 ;
        RECT 64.090 51.620 64.430 52.450 ;
        RECT 69.610 51.620 69.950 52.450 ;
        RECT 75.130 51.620 75.470 52.450 ;
        RECT 79.065 52.225 80.735 52.995 ;
        RECT 81.365 52.270 81.655 52.995 ;
        RECT 81.825 52.450 87.170 52.995 ;
        RECT 87.345 52.450 92.690 52.995 ;
        RECT 92.865 52.450 98.210 52.995 ;
        RECT 98.385 52.450 103.730 52.995 ;
        RECT 79.065 51.705 79.815 52.225 ;
        RECT 83.410 51.620 83.750 52.450 ;
        RECT 88.930 51.620 89.270 52.450 ;
        RECT 94.450 51.620 94.790 52.450 ;
        RECT 99.970 51.620 100.310 52.450 ;
        RECT 103.905 52.225 106.495 52.995 ;
        RECT 107.125 52.270 107.415 52.995 ;
        RECT 107.585 52.450 112.930 52.995 ;
        RECT 113.105 52.450 118.450 52.995 ;
        RECT 118.625 52.450 123.970 52.995 ;
        RECT 124.145 52.450 129.490 52.995 ;
        RECT 103.905 51.705 105.115 52.225 ;
        RECT 109.170 51.620 109.510 52.450 ;
        RECT 114.690 51.620 115.030 52.450 ;
        RECT 120.210 51.620 120.550 52.450 ;
        RECT 125.730 51.620 126.070 52.450 ;
        RECT 129.665 52.225 132.255 52.995 ;
        RECT 132.885 52.270 133.175 52.995 ;
        RECT 133.345 52.450 138.690 52.995 ;
        RECT 129.665 51.705 130.875 52.225 ;
        RECT 134.930 51.620 135.270 52.450 ;
        RECT 138.865 52.225 142.375 52.995 ;
        RECT 143.005 52.245 144.215 52.995 ;
        RECT 138.865 51.705 140.515 52.225 ;
        RECT 143.695 51.705 144.215 52.245 ;
        RECT 55.605 48.475 56.125 49.015 ;
        RECT 55.605 47.725 56.815 48.475 ;
        RECT 58.570 48.270 58.910 49.100 ;
        RECT 64.090 48.270 64.430 49.100 ;
        RECT 56.985 47.725 62.330 48.270 ;
        RECT 62.505 47.725 67.850 48.270 ;
        RECT 68.485 47.725 68.775 48.450 ;
        RECT 70.530 48.270 70.870 49.100 ;
        RECT 76.050 48.270 76.390 49.100 ;
        RECT 81.570 48.270 81.910 49.100 ;
        RECT 87.090 48.270 87.430 49.100 ;
        RECT 91.025 48.495 92.235 49.015 ;
        RECT 68.945 47.725 74.290 48.270 ;
        RECT 74.465 47.725 79.810 48.270 ;
        RECT 79.985 47.725 85.330 48.270 ;
        RECT 85.505 47.725 90.850 48.270 ;
        RECT 91.025 47.725 93.615 48.495 ;
        RECT 94.245 47.725 94.535 48.450 ;
        RECT 96.290 48.270 96.630 49.100 ;
        RECT 101.810 48.270 102.150 49.100 ;
        RECT 107.330 48.270 107.670 49.100 ;
        RECT 112.850 48.270 113.190 49.100 ;
        RECT 116.785 48.495 117.995 49.015 ;
        RECT 94.705 47.725 100.050 48.270 ;
        RECT 100.225 47.725 105.570 48.270 ;
        RECT 105.745 47.725 111.090 48.270 ;
        RECT 111.265 47.725 116.610 48.270 ;
        RECT 116.785 47.725 119.375 48.495 ;
        RECT 120.005 47.725 120.295 48.450 ;
        RECT 122.050 48.270 122.390 49.100 ;
        RECT 127.570 48.270 127.910 49.100 ;
        RECT 133.090 48.270 133.430 49.100 ;
        RECT 138.610 48.270 138.950 49.100 ;
        RECT 143.695 48.475 144.215 49.015 ;
        RECT 120.465 47.725 125.810 48.270 ;
        RECT 125.985 47.725 131.330 48.270 ;
        RECT 131.505 47.725 136.850 48.270 ;
        RECT 137.025 47.725 142.370 48.270 ;
        RECT 143.005 47.725 144.215 48.475 ;
        RECT 55.520 47.555 144.300 47.725 ;
        RECT 55.605 46.805 56.815 47.555 ;
        RECT 56.985 47.010 62.330 47.555 ;
        RECT 62.505 47.010 67.850 47.555 ;
        RECT 68.025 47.010 73.370 47.555 ;
        RECT 73.545 47.010 78.890 47.555 ;
        RECT 55.605 46.265 56.125 46.805 ;
        RECT 58.570 46.180 58.910 47.010 ;
        RECT 64.090 46.180 64.430 47.010 ;
        RECT 69.610 46.180 69.950 47.010 ;
        RECT 75.130 46.180 75.470 47.010 ;
        RECT 79.065 46.785 80.735 47.555 ;
        RECT 81.365 46.830 81.655 47.555 ;
        RECT 81.825 47.010 87.170 47.555 ;
        RECT 87.345 47.010 92.690 47.555 ;
        RECT 92.865 47.010 98.210 47.555 ;
        RECT 98.385 47.010 103.730 47.555 ;
        RECT 79.065 46.265 79.815 46.785 ;
        RECT 83.410 46.180 83.750 47.010 ;
        RECT 88.930 46.180 89.270 47.010 ;
        RECT 94.450 46.180 94.790 47.010 ;
        RECT 99.970 46.180 100.310 47.010 ;
        RECT 103.905 46.785 106.495 47.555 ;
        RECT 107.125 46.830 107.415 47.555 ;
        RECT 107.585 47.010 112.930 47.555 ;
        RECT 113.105 47.010 118.450 47.555 ;
        RECT 118.625 47.010 123.970 47.555 ;
        RECT 124.145 47.010 129.490 47.555 ;
        RECT 103.905 46.265 105.115 46.785 ;
        RECT 109.170 46.180 109.510 47.010 ;
        RECT 114.690 46.180 115.030 47.010 ;
        RECT 120.210 46.180 120.550 47.010 ;
        RECT 125.730 46.180 126.070 47.010 ;
        RECT 129.665 46.785 132.255 47.555 ;
        RECT 132.885 46.830 133.175 47.555 ;
        RECT 133.345 47.010 138.690 47.555 ;
        RECT 129.665 46.265 130.875 46.785 ;
        RECT 134.930 46.180 135.270 47.010 ;
        RECT 138.865 46.785 142.375 47.555 ;
        RECT 143.005 46.805 144.215 47.555 ;
        RECT 138.865 46.265 140.515 46.785 ;
        RECT 143.695 46.265 144.215 46.805 ;
        RECT 55.605 43.035 56.125 43.575 ;
        RECT 55.605 42.285 56.815 43.035 ;
        RECT 58.570 42.830 58.910 43.660 ;
        RECT 64.090 42.830 64.430 43.660 ;
        RECT 56.985 42.285 62.330 42.830 ;
        RECT 62.505 42.285 67.850 42.830 ;
        RECT 68.485 42.285 68.775 43.010 ;
        RECT 70.530 42.830 70.870 43.660 ;
        RECT 76.050 42.830 76.390 43.660 ;
        RECT 81.570 42.830 81.910 43.660 ;
        RECT 87.090 42.830 87.430 43.660 ;
        RECT 91.025 43.055 92.235 43.575 ;
        RECT 68.945 42.285 74.290 42.830 ;
        RECT 74.465 42.285 79.810 42.830 ;
        RECT 79.985 42.285 85.330 42.830 ;
        RECT 85.505 42.285 90.850 42.830 ;
        RECT 91.025 42.285 93.615 43.055 ;
        RECT 94.245 42.285 94.535 43.010 ;
        RECT 96.290 42.830 96.630 43.660 ;
        RECT 101.810 42.830 102.150 43.660 ;
        RECT 107.330 42.830 107.670 43.660 ;
        RECT 112.850 42.830 113.190 43.660 ;
        RECT 116.785 43.055 117.995 43.575 ;
        RECT 94.705 42.285 100.050 42.830 ;
        RECT 100.225 42.285 105.570 42.830 ;
        RECT 105.745 42.285 111.090 42.830 ;
        RECT 111.265 42.285 116.610 42.830 ;
        RECT 116.785 42.285 119.375 43.055 ;
        RECT 120.005 42.285 120.295 43.010 ;
        RECT 122.050 42.830 122.390 43.660 ;
        RECT 127.570 42.830 127.910 43.660 ;
        RECT 133.090 42.830 133.430 43.660 ;
        RECT 138.610 42.830 138.950 43.660 ;
        RECT 143.695 43.035 144.215 43.575 ;
        RECT 120.465 42.285 125.810 42.830 ;
        RECT 125.985 42.285 131.330 42.830 ;
        RECT 131.505 42.285 136.850 42.830 ;
        RECT 137.025 42.285 142.370 42.830 ;
        RECT 143.005 42.285 144.215 43.035 ;
        RECT 55.520 42.115 144.300 42.285 ;
        RECT 55.605 41.365 56.815 42.115 ;
        RECT 56.985 41.570 62.330 42.115 ;
        RECT 62.505 41.570 67.850 42.115 ;
        RECT 68.025 41.570 73.370 42.115 ;
        RECT 73.545 41.570 78.890 42.115 ;
        RECT 55.605 40.825 56.125 41.365 ;
        RECT 58.570 40.740 58.910 41.570 ;
        RECT 64.090 40.740 64.430 41.570 ;
        RECT 69.610 40.740 69.950 41.570 ;
        RECT 75.130 40.740 75.470 41.570 ;
        RECT 79.065 41.345 80.735 42.115 ;
        RECT 81.365 41.390 81.655 42.115 ;
        RECT 81.825 41.570 87.170 42.115 ;
        RECT 87.345 41.570 92.690 42.115 ;
        RECT 92.865 41.570 98.210 42.115 ;
        RECT 98.385 41.570 103.730 42.115 ;
        RECT 79.065 40.825 79.815 41.345 ;
        RECT 83.410 40.740 83.750 41.570 ;
        RECT 88.930 40.740 89.270 41.570 ;
        RECT 94.450 40.740 94.790 41.570 ;
        RECT 99.970 40.740 100.310 41.570 ;
        RECT 103.905 41.345 106.495 42.115 ;
        RECT 107.125 41.390 107.415 42.115 ;
        RECT 107.585 41.570 112.930 42.115 ;
        RECT 113.105 41.570 118.450 42.115 ;
        RECT 118.625 41.570 123.970 42.115 ;
        RECT 124.145 41.570 129.490 42.115 ;
        RECT 103.905 40.825 105.115 41.345 ;
        RECT 109.170 40.740 109.510 41.570 ;
        RECT 114.690 40.740 115.030 41.570 ;
        RECT 120.210 40.740 120.550 41.570 ;
        RECT 125.730 40.740 126.070 41.570 ;
        RECT 129.665 41.345 132.255 42.115 ;
        RECT 132.885 41.390 133.175 42.115 ;
        RECT 133.345 41.570 138.690 42.115 ;
        RECT 129.665 40.825 130.875 41.345 ;
        RECT 134.930 40.740 135.270 41.570 ;
        RECT 138.865 41.345 142.375 42.115 ;
        RECT 143.005 41.365 144.215 42.115 ;
        RECT 138.865 40.825 140.515 41.345 ;
        RECT 143.695 40.825 144.215 41.365 ;
        RECT 55.605 37.595 56.125 38.135 ;
        RECT 55.605 36.845 56.815 37.595 ;
        RECT 58.570 37.390 58.910 38.220 ;
        RECT 64.090 37.390 64.430 38.220 ;
        RECT 56.985 36.845 62.330 37.390 ;
        RECT 62.505 36.845 67.850 37.390 ;
        RECT 68.485 36.845 68.775 37.570 ;
        RECT 70.530 37.390 70.870 38.220 ;
        RECT 76.050 37.390 76.390 38.220 ;
        RECT 81.570 37.390 81.910 38.220 ;
        RECT 87.090 37.390 87.430 38.220 ;
        RECT 91.025 37.615 92.235 38.135 ;
        RECT 68.945 36.845 74.290 37.390 ;
        RECT 74.465 36.845 79.810 37.390 ;
        RECT 79.985 36.845 85.330 37.390 ;
        RECT 85.505 36.845 90.850 37.390 ;
        RECT 91.025 36.845 93.615 37.615 ;
        RECT 94.245 36.845 94.535 37.570 ;
        RECT 96.290 37.390 96.630 38.220 ;
        RECT 101.810 37.390 102.150 38.220 ;
        RECT 107.330 37.390 107.670 38.220 ;
        RECT 112.850 37.390 113.190 38.220 ;
        RECT 116.785 37.615 117.995 38.135 ;
        RECT 94.705 36.845 100.050 37.390 ;
        RECT 100.225 36.845 105.570 37.390 ;
        RECT 105.745 36.845 111.090 37.390 ;
        RECT 111.265 36.845 116.610 37.390 ;
        RECT 116.785 36.845 119.375 37.615 ;
        RECT 120.005 36.845 120.295 37.570 ;
        RECT 122.050 37.390 122.390 38.220 ;
        RECT 127.570 37.390 127.910 38.220 ;
        RECT 133.090 37.390 133.430 38.220 ;
        RECT 138.610 37.390 138.950 38.220 ;
        RECT 143.695 37.595 144.215 38.135 ;
        RECT 120.465 36.845 125.810 37.390 ;
        RECT 125.985 36.845 131.330 37.390 ;
        RECT 131.505 36.845 136.850 37.390 ;
        RECT 137.025 36.845 142.370 37.390 ;
        RECT 143.005 36.845 144.215 37.595 ;
        RECT 55.520 36.675 144.300 36.845 ;
        RECT 55.605 35.925 56.815 36.675 ;
        RECT 56.985 36.130 62.330 36.675 ;
        RECT 62.505 36.130 67.850 36.675 ;
        RECT 68.025 36.130 73.370 36.675 ;
        RECT 73.545 36.130 78.890 36.675 ;
        RECT 55.605 35.385 56.125 35.925 ;
        RECT 58.570 35.300 58.910 36.130 ;
        RECT 64.090 35.300 64.430 36.130 ;
        RECT 69.610 35.300 69.950 36.130 ;
        RECT 75.130 35.300 75.470 36.130 ;
        RECT 79.065 35.905 80.735 36.675 ;
        RECT 81.365 35.950 81.655 36.675 ;
        RECT 81.825 36.130 87.170 36.675 ;
        RECT 87.345 36.130 92.690 36.675 ;
        RECT 92.865 36.130 98.210 36.675 ;
        RECT 98.385 36.130 103.730 36.675 ;
        RECT 79.065 35.385 79.815 35.905 ;
        RECT 83.410 35.300 83.750 36.130 ;
        RECT 88.930 35.300 89.270 36.130 ;
        RECT 94.450 35.300 94.790 36.130 ;
        RECT 99.970 35.300 100.310 36.130 ;
        RECT 103.905 35.905 106.495 36.675 ;
        RECT 107.125 35.950 107.415 36.675 ;
        RECT 107.585 36.130 112.930 36.675 ;
        RECT 113.105 36.130 118.450 36.675 ;
        RECT 118.625 36.130 123.970 36.675 ;
        RECT 124.145 36.130 129.490 36.675 ;
        RECT 103.905 35.385 105.115 35.905 ;
        RECT 109.170 35.300 109.510 36.130 ;
        RECT 114.690 35.300 115.030 36.130 ;
        RECT 120.210 35.300 120.550 36.130 ;
        RECT 125.730 35.300 126.070 36.130 ;
        RECT 129.665 35.905 132.255 36.675 ;
        RECT 132.885 35.950 133.175 36.675 ;
        RECT 133.345 36.130 138.690 36.675 ;
        RECT 129.665 35.385 130.875 35.905 ;
        RECT 134.930 35.300 135.270 36.130 ;
        RECT 138.865 35.905 142.375 36.675 ;
        RECT 143.005 35.925 144.215 36.675 ;
        RECT 138.865 35.385 140.515 35.905 ;
        RECT 143.695 35.385 144.215 35.925 ;
        RECT 55.605 32.155 56.125 32.695 ;
        RECT 55.605 31.405 56.815 32.155 ;
        RECT 58.570 31.950 58.910 32.780 ;
        RECT 64.090 31.950 64.430 32.780 ;
        RECT 56.985 31.405 62.330 31.950 ;
        RECT 62.505 31.405 67.850 31.950 ;
        RECT 68.485 31.405 68.775 32.130 ;
        RECT 70.530 31.950 70.870 32.780 ;
        RECT 76.050 31.950 76.390 32.780 ;
        RECT 81.570 31.950 81.910 32.780 ;
        RECT 87.090 31.950 87.430 32.780 ;
        RECT 91.025 32.175 92.235 32.695 ;
        RECT 68.945 31.405 74.290 31.950 ;
        RECT 74.465 31.405 79.810 31.950 ;
        RECT 79.985 31.405 85.330 31.950 ;
        RECT 85.505 31.405 90.850 31.950 ;
        RECT 91.025 31.405 93.615 32.175 ;
        RECT 94.245 31.405 94.535 32.130 ;
        RECT 96.290 31.950 96.630 32.780 ;
        RECT 101.810 31.950 102.150 32.780 ;
        RECT 107.330 31.950 107.670 32.780 ;
        RECT 112.850 31.950 113.190 32.780 ;
        RECT 116.785 32.175 117.995 32.695 ;
        RECT 94.705 31.405 100.050 31.950 ;
        RECT 100.225 31.405 105.570 31.950 ;
        RECT 105.745 31.405 111.090 31.950 ;
        RECT 111.265 31.405 116.610 31.950 ;
        RECT 116.785 31.405 119.375 32.175 ;
        RECT 120.005 31.405 120.295 32.130 ;
        RECT 122.050 31.950 122.390 32.780 ;
        RECT 127.570 31.950 127.910 32.780 ;
        RECT 133.090 31.950 133.430 32.780 ;
        RECT 138.610 31.950 138.950 32.780 ;
        RECT 143.695 32.155 144.215 32.695 ;
        RECT 120.465 31.405 125.810 31.950 ;
        RECT 125.985 31.405 131.330 31.950 ;
        RECT 131.505 31.405 136.850 31.950 ;
        RECT 137.025 31.405 142.370 31.950 ;
        RECT 143.005 31.405 144.215 32.155 ;
        RECT 55.520 31.235 144.300 31.405 ;
        RECT 55.605 30.485 56.815 31.235 ;
        RECT 56.985 30.690 62.330 31.235 ;
        RECT 62.505 30.690 67.850 31.235 ;
        RECT 68.025 30.690 73.370 31.235 ;
        RECT 73.545 30.690 78.890 31.235 ;
        RECT 55.605 29.945 56.125 30.485 ;
        RECT 58.570 29.860 58.910 30.690 ;
        RECT 64.090 29.860 64.430 30.690 ;
        RECT 69.610 29.860 69.950 30.690 ;
        RECT 75.130 29.860 75.470 30.690 ;
        RECT 79.065 30.465 80.735 31.235 ;
        RECT 81.365 30.510 81.655 31.235 ;
        RECT 81.825 30.690 87.170 31.235 ;
        RECT 87.345 30.690 92.690 31.235 ;
        RECT 92.865 30.690 98.210 31.235 ;
        RECT 98.385 30.690 103.730 31.235 ;
        RECT 79.065 29.945 79.815 30.465 ;
        RECT 83.410 29.860 83.750 30.690 ;
        RECT 88.930 29.860 89.270 30.690 ;
        RECT 94.450 29.860 94.790 30.690 ;
        RECT 99.970 29.860 100.310 30.690 ;
        RECT 103.905 30.465 106.495 31.235 ;
        RECT 107.125 30.510 107.415 31.235 ;
        RECT 107.585 30.690 112.930 31.235 ;
        RECT 113.105 30.690 118.450 31.235 ;
        RECT 118.625 30.690 123.970 31.235 ;
        RECT 124.145 30.690 129.490 31.235 ;
        RECT 103.905 29.945 105.115 30.465 ;
        RECT 109.170 29.860 109.510 30.690 ;
        RECT 114.690 29.860 115.030 30.690 ;
        RECT 120.210 29.860 120.550 30.690 ;
        RECT 125.730 29.860 126.070 30.690 ;
        RECT 129.665 30.465 132.255 31.235 ;
        RECT 132.885 30.510 133.175 31.235 ;
        RECT 133.345 30.690 138.690 31.235 ;
        RECT 129.665 29.945 130.875 30.465 ;
        RECT 134.930 29.860 135.270 30.690 ;
        RECT 138.865 30.465 142.375 31.235 ;
        RECT 143.005 30.485 144.215 31.235 ;
        RECT 138.865 29.945 140.515 30.465 ;
        RECT 143.695 29.945 144.215 30.485 ;
        RECT 55.605 26.715 56.125 27.255 ;
        RECT 55.605 25.965 56.815 26.715 ;
        RECT 58.570 26.510 58.910 27.340 ;
        RECT 64.090 26.510 64.430 27.340 ;
        RECT 56.985 25.965 62.330 26.510 ;
        RECT 62.505 25.965 67.850 26.510 ;
        RECT 68.485 25.965 68.775 26.690 ;
        RECT 70.530 26.510 70.870 27.340 ;
        RECT 76.050 26.510 76.390 27.340 ;
        RECT 79.985 26.715 80.505 27.255 ;
        RECT 68.945 25.965 74.290 26.510 ;
        RECT 74.465 25.965 79.810 26.510 ;
        RECT 79.985 25.965 81.195 26.715 ;
        RECT 81.365 25.965 81.655 26.690 ;
        RECT 83.410 26.510 83.750 27.340 ;
        RECT 88.930 26.510 89.270 27.340 ;
        RECT 92.865 26.715 93.385 27.255 ;
        RECT 81.825 25.965 87.170 26.510 ;
        RECT 87.345 25.965 92.690 26.510 ;
        RECT 92.865 25.965 94.075 26.715 ;
        RECT 94.245 25.965 94.535 26.690 ;
        RECT 96.290 26.510 96.630 27.340 ;
        RECT 101.810 26.510 102.150 27.340 ;
        RECT 105.745 26.715 106.265 27.255 ;
        RECT 94.705 25.965 100.050 26.510 ;
        RECT 100.225 25.965 105.570 26.510 ;
        RECT 105.745 25.965 106.955 26.715 ;
        RECT 107.125 25.965 107.415 26.690 ;
        RECT 109.170 26.510 109.510 27.340 ;
        RECT 114.690 26.510 115.030 27.340 ;
        RECT 118.625 26.715 119.145 27.255 ;
        RECT 107.585 25.965 112.930 26.510 ;
        RECT 113.105 25.965 118.450 26.510 ;
        RECT 118.625 25.965 119.835 26.715 ;
        RECT 120.005 25.965 120.295 26.690 ;
        RECT 122.050 26.510 122.390 27.340 ;
        RECT 127.570 26.510 127.910 27.340 ;
        RECT 131.505 26.715 132.025 27.255 ;
        RECT 120.465 25.965 125.810 26.510 ;
        RECT 125.985 25.965 131.330 26.510 ;
        RECT 131.505 25.965 132.715 26.715 ;
        RECT 132.885 25.965 133.175 26.690 ;
        RECT 134.930 26.510 135.270 27.340 ;
        RECT 138.865 26.735 140.515 27.255 ;
        RECT 133.345 25.965 138.690 26.510 ;
        RECT 138.865 25.965 142.375 26.735 ;
        RECT 143.695 26.715 144.215 27.255 ;
        RECT 143.005 25.965 144.215 26.715 ;
        RECT 55.520 25.795 144.300 25.965 ;
      LAYER mcon ;
        RECT 55.665 101.955 55.835 102.125 ;
        RECT 56.125 101.955 56.295 102.125 ;
        RECT 56.585 101.955 56.755 102.125 ;
        RECT 57.045 101.955 57.215 102.125 ;
        RECT 57.505 101.955 57.675 102.125 ;
        RECT 57.965 101.955 58.135 102.125 ;
        RECT 58.425 101.955 58.595 102.125 ;
        RECT 58.885 101.955 59.055 102.125 ;
        RECT 59.345 101.955 59.515 102.125 ;
        RECT 59.805 101.955 59.975 102.125 ;
        RECT 60.265 101.955 60.435 102.125 ;
        RECT 60.725 101.955 60.895 102.125 ;
        RECT 61.185 101.955 61.355 102.125 ;
        RECT 61.645 101.955 61.815 102.125 ;
        RECT 62.105 101.955 62.275 102.125 ;
        RECT 62.565 101.955 62.735 102.125 ;
        RECT 63.025 101.955 63.195 102.125 ;
        RECT 63.485 101.955 63.655 102.125 ;
        RECT 63.945 101.955 64.115 102.125 ;
        RECT 64.405 101.955 64.575 102.125 ;
        RECT 64.865 101.955 65.035 102.125 ;
        RECT 65.325 101.955 65.495 102.125 ;
        RECT 65.785 101.955 65.955 102.125 ;
        RECT 66.245 101.955 66.415 102.125 ;
        RECT 66.705 101.955 66.875 102.125 ;
        RECT 67.165 101.955 67.335 102.125 ;
        RECT 67.625 101.955 67.795 102.125 ;
        RECT 68.085 101.955 68.255 102.125 ;
        RECT 68.545 101.955 68.715 102.125 ;
        RECT 69.005 101.955 69.175 102.125 ;
        RECT 69.465 101.955 69.635 102.125 ;
        RECT 69.925 101.955 70.095 102.125 ;
        RECT 70.385 101.955 70.555 102.125 ;
        RECT 70.845 101.955 71.015 102.125 ;
        RECT 71.305 101.955 71.475 102.125 ;
        RECT 71.765 101.955 71.935 102.125 ;
        RECT 72.225 101.955 72.395 102.125 ;
        RECT 72.685 101.955 72.855 102.125 ;
        RECT 73.145 101.955 73.315 102.125 ;
        RECT 73.605 101.955 73.775 102.125 ;
        RECT 74.065 101.955 74.235 102.125 ;
        RECT 74.525 101.955 74.695 102.125 ;
        RECT 74.985 101.955 75.155 102.125 ;
        RECT 75.445 101.955 75.615 102.125 ;
        RECT 75.905 101.955 76.075 102.125 ;
        RECT 76.365 101.955 76.535 102.125 ;
        RECT 76.825 101.955 76.995 102.125 ;
        RECT 77.285 101.955 77.455 102.125 ;
        RECT 77.745 101.955 77.915 102.125 ;
        RECT 78.205 101.955 78.375 102.125 ;
        RECT 78.665 101.955 78.835 102.125 ;
        RECT 79.125 101.955 79.295 102.125 ;
        RECT 79.585 101.955 79.755 102.125 ;
        RECT 80.045 101.955 80.215 102.125 ;
        RECT 80.505 101.955 80.675 102.125 ;
        RECT 80.965 101.955 81.135 102.125 ;
        RECT 81.425 101.955 81.595 102.125 ;
        RECT 81.885 101.955 82.055 102.125 ;
        RECT 82.345 101.955 82.515 102.125 ;
        RECT 82.805 101.955 82.975 102.125 ;
        RECT 83.265 101.955 83.435 102.125 ;
        RECT 83.725 101.955 83.895 102.125 ;
        RECT 84.185 101.955 84.355 102.125 ;
        RECT 84.645 101.955 84.815 102.125 ;
        RECT 85.105 101.955 85.275 102.125 ;
        RECT 85.565 101.955 85.735 102.125 ;
        RECT 86.025 101.955 86.195 102.125 ;
        RECT 86.485 101.955 86.655 102.125 ;
        RECT 86.945 101.955 87.115 102.125 ;
        RECT 87.405 101.955 87.575 102.125 ;
        RECT 87.865 101.955 88.035 102.125 ;
        RECT 88.325 101.955 88.495 102.125 ;
        RECT 88.785 101.955 88.955 102.125 ;
        RECT 89.245 101.955 89.415 102.125 ;
        RECT 89.705 101.955 89.875 102.125 ;
        RECT 90.165 101.955 90.335 102.125 ;
        RECT 90.625 101.955 90.795 102.125 ;
        RECT 91.085 101.955 91.255 102.125 ;
        RECT 91.545 101.955 91.715 102.125 ;
        RECT 92.005 101.955 92.175 102.125 ;
        RECT 92.465 101.955 92.635 102.125 ;
        RECT 92.925 101.955 93.095 102.125 ;
        RECT 93.385 101.955 93.555 102.125 ;
        RECT 93.845 101.955 94.015 102.125 ;
        RECT 94.305 101.955 94.475 102.125 ;
        RECT 94.765 101.955 94.935 102.125 ;
        RECT 95.225 101.955 95.395 102.125 ;
        RECT 95.685 101.955 95.855 102.125 ;
        RECT 96.145 101.955 96.315 102.125 ;
        RECT 96.605 101.955 96.775 102.125 ;
        RECT 97.065 101.955 97.235 102.125 ;
        RECT 97.525 101.955 97.695 102.125 ;
        RECT 97.985 101.955 98.155 102.125 ;
        RECT 98.445 101.955 98.615 102.125 ;
        RECT 98.905 101.955 99.075 102.125 ;
        RECT 99.365 101.955 99.535 102.125 ;
        RECT 99.825 101.955 99.995 102.125 ;
        RECT 100.285 101.955 100.455 102.125 ;
        RECT 100.745 101.955 100.915 102.125 ;
        RECT 101.205 101.955 101.375 102.125 ;
        RECT 101.665 101.955 101.835 102.125 ;
        RECT 102.125 101.955 102.295 102.125 ;
        RECT 102.585 101.955 102.755 102.125 ;
        RECT 103.045 101.955 103.215 102.125 ;
        RECT 103.505 101.955 103.675 102.125 ;
        RECT 103.965 101.955 104.135 102.125 ;
        RECT 104.425 101.955 104.595 102.125 ;
        RECT 104.885 101.955 105.055 102.125 ;
        RECT 105.345 101.955 105.515 102.125 ;
        RECT 105.805 101.955 105.975 102.125 ;
        RECT 106.265 101.955 106.435 102.125 ;
        RECT 106.725 101.955 106.895 102.125 ;
        RECT 107.185 101.955 107.355 102.125 ;
        RECT 107.645 101.955 107.815 102.125 ;
        RECT 108.105 101.955 108.275 102.125 ;
        RECT 108.565 101.955 108.735 102.125 ;
        RECT 109.025 101.955 109.195 102.125 ;
        RECT 109.485 101.955 109.655 102.125 ;
        RECT 109.945 101.955 110.115 102.125 ;
        RECT 110.405 101.955 110.575 102.125 ;
        RECT 110.865 101.955 111.035 102.125 ;
        RECT 111.325 101.955 111.495 102.125 ;
        RECT 111.785 101.955 111.955 102.125 ;
        RECT 112.245 101.955 112.415 102.125 ;
        RECT 112.705 101.955 112.875 102.125 ;
        RECT 113.165 101.955 113.335 102.125 ;
        RECT 113.625 101.955 113.795 102.125 ;
        RECT 114.085 101.955 114.255 102.125 ;
        RECT 114.545 101.955 114.715 102.125 ;
        RECT 115.005 101.955 115.175 102.125 ;
        RECT 115.465 101.955 115.635 102.125 ;
        RECT 115.925 101.955 116.095 102.125 ;
        RECT 116.385 101.955 116.555 102.125 ;
        RECT 116.845 101.955 117.015 102.125 ;
        RECT 117.305 101.955 117.475 102.125 ;
        RECT 117.765 101.955 117.935 102.125 ;
        RECT 118.225 101.955 118.395 102.125 ;
        RECT 118.685 101.955 118.855 102.125 ;
        RECT 119.145 101.955 119.315 102.125 ;
        RECT 119.605 101.955 119.775 102.125 ;
        RECT 120.065 101.955 120.235 102.125 ;
        RECT 120.525 101.955 120.695 102.125 ;
        RECT 120.985 101.955 121.155 102.125 ;
        RECT 121.445 101.955 121.615 102.125 ;
        RECT 121.905 101.955 122.075 102.125 ;
        RECT 122.365 101.955 122.535 102.125 ;
        RECT 122.825 101.955 122.995 102.125 ;
        RECT 123.285 101.955 123.455 102.125 ;
        RECT 123.745 101.955 123.915 102.125 ;
        RECT 124.205 101.955 124.375 102.125 ;
        RECT 124.665 101.955 124.835 102.125 ;
        RECT 125.125 101.955 125.295 102.125 ;
        RECT 125.585 101.955 125.755 102.125 ;
        RECT 126.045 101.955 126.215 102.125 ;
        RECT 126.505 101.955 126.675 102.125 ;
        RECT 126.965 101.955 127.135 102.125 ;
        RECT 127.425 101.955 127.595 102.125 ;
        RECT 127.885 101.955 128.055 102.125 ;
        RECT 128.345 101.955 128.515 102.125 ;
        RECT 128.805 101.955 128.975 102.125 ;
        RECT 129.265 101.955 129.435 102.125 ;
        RECT 129.725 101.955 129.895 102.125 ;
        RECT 130.185 101.955 130.355 102.125 ;
        RECT 130.645 101.955 130.815 102.125 ;
        RECT 131.105 101.955 131.275 102.125 ;
        RECT 131.565 101.955 131.735 102.125 ;
        RECT 132.025 101.955 132.195 102.125 ;
        RECT 132.485 101.955 132.655 102.125 ;
        RECT 132.945 101.955 133.115 102.125 ;
        RECT 133.405 101.955 133.575 102.125 ;
        RECT 133.865 101.955 134.035 102.125 ;
        RECT 134.325 101.955 134.495 102.125 ;
        RECT 134.785 101.955 134.955 102.125 ;
        RECT 135.245 101.955 135.415 102.125 ;
        RECT 135.705 101.955 135.875 102.125 ;
        RECT 136.165 101.955 136.335 102.125 ;
        RECT 136.625 101.955 136.795 102.125 ;
        RECT 137.085 101.955 137.255 102.125 ;
        RECT 137.545 101.955 137.715 102.125 ;
        RECT 138.005 101.955 138.175 102.125 ;
        RECT 138.465 101.955 138.635 102.125 ;
        RECT 138.925 101.955 139.095 102.125 ;
        RECT 139.385 101.955 139.555 102.125 ;
        RECT 139.845 101.955 140.015 102.125 ;
        RECT 140.305 101.955 140.475 102.125 ;
        RECT 140.765 101.955 140.935 102.125 ;
        RECT 141.225 101.955 141.395 102.125 ;
        RECT 141.685 101.955 141.855 102.125 ;
        RECT 142.145 101.955 142.315 102.125 ;
        RECT 142.605 101.955 142.775 102.125 ;
        RECT 143.065 101.955 143.235 102.125 ;
        RECT 143.525 101.955 143.695 102.125 ;
        RECT 143.985 101.955 144.155 102.125 ;
        RECT 55.665 96.515 55.835 96.685 ;
        RECT 56.125 96.515 56.295 96.685 ;
        RECT 56.585 96.515 56.755 96.685 ;
        RECT 57.045 96.515 57.215 96.685 ;
        RECT 57.505 96.515 57.675 96.685 ;
        RECT 57.965 96.515 58.135 96.685 ;
        RECT 58.425 96.515 58.595 96.685 ;
        RECT 58.885 96.515 59.055 96.685 ;
        RECT 59.345 96.515 59.515 96.685 ;
        RECT 59.805 96.515 59.975 96.685 ;
        RECT 60.265 96.515 60.435 96.685 ;
        RECT 60.725 96.515 60.895 96.685 ;
        RECT 61.185 96.515 61.355 96.685 ;
        RECT 61.645 96.515 61.815 96.685 ;
        RECT 62.105 96.515 62.275 96.685 ;
        RECT 62.565 96.515 62.735 96.685 ;
        RECT 63.025 96.515 63.195 96.685 ;
        RECT 63.485 96.515 63.655 96.685 ;
        RECT 63.945 96.515 64.115 96.685 ;
        RECT 64.405 96.515 64.575 96.685 ;
        RECT 64.865 96.515 65.035 96.685 ;
        RECT 65.325 96.515 65.495 96.685 ;
        RECT 65.785 96.515 65.955 96.685 ;
        RECT 66.245 96.515 66.415 96.685 ;
        RECT 66.705 96.515 66.875 96.685 ;
        RECT 67.165 96.515 67.335 96.685 ;
        RECT 67.625 96.515 67.795 96.685 ;
        RECT 68.085 96.515 68.255 96.685 ;
        RECT 68.545 96.515 68.715 96.685 ;
        RECT 69.005 96.515 69.175 96.685 ;
        RECT 69.465 96.515 69.635 96.685 ;
        RECT 69.925 96.515 70.095 96.685 ;
        RECT 70.385 96.515 70.555 96.685 ;
        RECT 70.845 96.515 71.015 96.685 ;
        RECT 71.305 96.515 71.475 96.685 ;
        RECT 71.765 96.515 71.935 96.685 ;
        RECT 72.225 96.515 72.395 96.685 ;
        RECT 72.685 96.515 72.855 96.685 ;
        RECT 73.145 96.515 73.315 96.685 ;
        RECT 73.605 96.515 73.775 96.685 ;
        RECT 74.065 96.515 74.235 96.685 ;
        RECT 74.525 96.515 74.695 96.685 ;
        RECT 74.985 96.515 75.155 96.685 ;
        RECT 75.445 96.515 75.615 96.685 ;
        RECT 75.905 96.515 76.075 96.685 ;
        RECT 76.365 96.515 76.535 96.685 ;
        RECT 76.825 96.515 76.995 96.685 ;
        RECT 77.285 96.515 77.455 96.685 ;
        RECT 77.745 96.515 77.915 96.685 ;
        RECT 78.205 96.515 78.375 96.685 ;
        RECT 78.665 96.515 78.835 96.685 ;
        RECT 79.125 96.515 79.295 96.685 ;
        RECT 79.585 96.515 79.755 96.685 ;
        RECT 80.045 96.515 80.215 96.685 ;
        RECT 80.505 96.515 80.675 96.685 ;
        RECT 80.965 96.515 81.135 96.685 ;
        RECT 81.425 96.515 81.595 96.685 ;
        RECT 81.885 96.515 82.055 96.685 ;
        RECT 82.345 96.515 82.515 96.685 ;
        RECT 82.805 96.515 82.975 96.685 ;
        RECT 83.265 96.515 83.435 96.685 ;
        RECT 83.725 96.515 83.895 96.685 ;
        RECT 84.185 96.515 84.355 96.685 ;
        RECT 84.645 96.515 84.815 96.685 ;
        RECT 85.105 96.515 85.275 96.685 ;
        RECT 85.565 96.515 85.735 96.685 ;
        RECT 86.025 96.515 86.195 96.685 ;
        RECT 86.485 96.515 86.655 96.685 ;
        RECT 86.945 96.515 87.115 96.685 ;
        RECT 87.405 96.515 87.575 96.685 ;
        RECT 87.865 96.515 88.035 96.685 ;
        RECT 88.325 96.515 88.495 96.685 ;
        RECT 88.785 96.515 88.955 96.685 ;
        RECT 89.245 96.515 89.415 96.685 ;
        RECT 89.705 96.515 89.875 96.685 ;
        RECT 90.165 96.515 90.335 96.685 ;
        RECT 90.625 96.515 90.795 96.685 ;
        RECT 91.085 96.515 91.255 96.685 ;
        RECT 91.545 96.515 91.715 96.685 ;
        RECT 92.005 96.515 92.175 96.685 ;
        RECT 92.465 96.515 92.635 96.685 ;
        RECT 92.925 96.515 93.095 96.685 ;
        RECT 93.385 96.515 93.555 96.685 ;
        RECT 93.845 96.515 94.015 96.685 ;
        RECT 94.305 96.515 94.475 96.685 ;
        RECT 94.765 96.515 94.935 96.685 ;
        RECT 95.225 96.515 95.395 96.685 ;
        RECT 95.685 96.515 95.855 96.685 ;
        RECT 96.145 96.515 96.315 96.685 ;
        RECT 96.605 96.515 96.775 96.685 ;
        RECT 97.065 96.515 97.235 96.685 ;
        RECT 97.525 96.515 97.695 96.685 ;
        RECT 97.985 96.515 98.155 96.685 ;
        RECT 98.445 96.515 98.615 96.685 ;
        RECT 98.905 96.515 99.075 96.685 ;
        RECT 99.365 96.515 99.535 96.685 ;
        RECT 99.825 96.515 99.995 96.685 ;
        RECT 100.285 96.515 100.455 96.685 ;
        RECT 100.745 96.515 100.915 96.685 ;
        RECT 101.205 96.515 101.375 96.685 ;
        RECT 101.665 96.515 101.835 96.685 ;
        RECT 102.125 96.515 102.295 96.685 ;
        RECT 102.585 96.515 102.755 96.685 ;
        RECT 103.045 96.515 103.215 96.685 ;
        RECT 103.505 96.515 103.675 96.685 ;
        RECT 103.965 96.515 104.135 96.685 ;
        RECT 104.425 96.515 104.595 96.685 ;
        RECT 104.885 96.515 105.055 96.685 ;
        RECT 105.345 96.515 105.515 96.685 ;
        RECT 105.805 96.515 105.975 96.685 ;
        RECT 106.265 96.515 106.435 96.685 ;
        RECT 106.725 96.515 106.895 96.685 ;
        RECT 107.185 96.515 107.355 96.685 ;
        RECT 107.645 96.515 107.815 96.685 ;
        RECT 108.105 96.515 108.275 96.685 ;
        RECT 108.565 96.515 108.735 96.685 ;
        RECT 109.025 96.515 109.195 96.685 ;
        RECT 109.485 96.515 109.655 96.685 ;
        RECT 109.945 96.515 110.115 96.685 ;
        RECT 110.405 96.515 110.575 96.685 ;
        RECT 110.865 96.515 111.035 96.685 ;
        RECT 111.325 96.515 111.495 96.685 ;
        RECT 111.785 96.515 111.955 96.685 ;
        RECT 112.245 96.515 112.415 96.685 ;
        RECT 112.705 96.515 112.875 96.685 ;
        RECT 113.165 96.515 113.335 96.685 ;
        RECT 113.625 96.515 113.795 96.685 ;
        RECT 114.085 96.515 114.255 96.685 ;
        RECT 114.545 96.515 114.715 96.685 ;
        RECT 115.005 96.515 115.175 96.685 ;
        RECT 115.465 96.515 115.635 96.685 ;
        RECT 115.925 96.515 116.095 96.685 ;
        RECT 116.385 96.515 116.555 96.685 ;
        RECT 116.845 96.515 117.015 96.685 ;
        RECT 117.305 96.515 117.475 96.685 ;
        RECT 117.765 96.515 117.935 96.685 ;
        RECT 118.225 96.515 118.395 96.685 ;
        RECT 118.685 96.515 118.855 96.685 ;
        RECT 119.145 96.515 119.315 96.685 ;
        RECT 119.605 96.515 119.775 96.685 ;
        RECT 120.065 96.515 120.235 96.685 ;
        RECT 120.525 96.515 120.695 96.685 ;
        RECT 120.985 96.515 121.155 96.685 ;
        RECT 121.445 96.515 121.615 96.685 ;
        RECT 121.905 96.515 122.075 96.685 ;
        RECT 122.365 96.515 122.535 96.685 ;
        RECT 122.825 96.515 122.995 96.685 ;
        RECT 123.285 96.515 123.455 96.685 ;
        RECT 123.745 96.515 123.915 96.685 ;
        RECT 124.205 96.515 124.375 96.685 ;
        RECT 124.665 96.515 124.835 96.685 ;
        RECT 125.125 96.515 125.295 96.685 ;
        RECT 125.585 96.515 125.755 96.685 ;
        RECT 126.045 96.515 126.215 96.685 ;
        RECT 126.505 96.515 126.675 96.685 ;
        RECT 126.965 96.515 127.135 96.685 ;
        RECT 127.425 96.515 127.595 96.685 ;
        RECT 127.885 96.515 128.055 96.685 ;
        RECT 128.345 96.515 128.515 96.685 ;
        RECT 128.805 96.515 128.975 96.685 ;
        RECT 129.265 96.515 129.435 96.685 ;
        RECT 129.725 96.515 129.895 96.685 ;
        RECT 130.185 96.515 130.355 96.685 ;
        RECT 130.645 96.515 130.815 96.685 ;
        RECT 131.105 96.515 131.275 96.685 ;
        RECT 131.565 96.515 131.735 96.685 ;
        RECT 132.025 96.515 132.195 96.685 ;
        RECT 132.485 96.515 132.655 96.685 ;
        RECT 132.945 96.515 133.115 96.685 ;
        RECT 133.405 96.515 133.575 96.685 ;
        RECT 133.865 96.515 134.035 96.685 ;
        RECT 134.325 96.515 134.495 96.685 ;
        RECT 134.785 96.515 134.955 96.685 ;
        RECT 135.245 96.515 135.415 96.685 ;
        RECT 135.705 96.515 135.875 96.685 ;
        RECT 136.165 96.515 136.335 96.685 ;
        RECT 136.625 96.515 136.795 96.685 ;
        RECT 137.085 96.515 137.255 96.685 ;
        RECT 137.545 96.515 137.715 96.685 ;
        RECT 138.005 96.515 138.175 96.685 ;
        RECT 138.465 96.515 138.635 96.685 ;
        RECT 138.925 96.515 139.095 96.685 ;
        RECT 139.385 96.515 139.555 96.685 ;
        RECT 139.845 96.515 140.015 96.685 ;
        RECT 140.305 96.515 140.475 96.685 ;
        RECT 140.765 96.515 140.935 96.685 ;
        RECT 141.225 96.515 141.395 96.685 ;
        RECT 141.685 96.515 141.855 96.685 ;
        RECT 142.145 96.515 142.315 96.685 ;
        RECT 142.605 96.515 142.775 96.685 ;
        RECT 143.065 96.515 143.235 96.685 ;
        RECT 143.525 96.515 143.695 96.685 ;
        RECT 143.985 96.515 144.155 96.685 ;
        RECT 55.665 91.075 55.835 91.245 ;
        RECT 56.125 91.075 56.295 91.245 ;
        RECT 56.585 91.075 56.755 91.245 ;
        RECT 57.045 91.075 57.215 91.245 ;
        RECT 57.505 91.075 57.675 91.245 ;
        RECT 57.965 91.075 58.135 91.245 ;
        RECT 58.425 91.075 58.595 91.245 ;
        RECT 58.885 91.075 59.055 91.245 ;
        RECT 59.345 91.075 59.515 91.245 ;
        RECT 59.805 91.075 59.975 91.245 ;
        RECT 60.265 91.075 60.435 91.245 ;
        RECT 60.725 91.075 60.895 91.245 ;
        RECT 61.185 91.075 61.355 91.245 ;
        RECT 61.645 91.075 61.815 91.245 ;
        RECT 62.105 91.075 62.275 91.245 ;
        RECT 62.565 91.075 62.735 91.245 ;
        RECT 63.025 91.075 63.195 91.245 ;
        RECT 63.485 91.075 63.655 91.245 ;
        RECT 63.945 91.075 64.115 91.245 ;
        RECT 64.405 91.075 64.575 91.245 ;
        RECT 64.865 91.075 65.035 91.245 ;
        RECT 65.325 91.075 65.495 91.245 ;
        RECT 65.785 91.075 65.955 91.245 ;
        RECT 66.245 91.075 66.415 91.245 ;
        RECT 66.705 91.075 66.875 91.245 ;
        RECT 67.165 91.075 67.335 91.245 ;
        RECT 67.625 91.075 67.795 91.245 ;
        RECT 68.085 91.075 68.255 91.245 ;
        RECT 68.545 91.075 68.715 91.245 ;
        RECT 69.005 91.075 69.175 91.245 ;
        RECT 69.465 91.075 69.635 91.245 ;
        RECT 69.925 91.075 70.095 91.245 ;
        RECT 70.385 91.075 70.555 91.245 ;
        RECT 70.845 91.075 71.015 91.245 ;
        RECT 71.305 91.075 71.475 91.245 ;
        RECT 71.765 91.075 71.935 91.245 ;
        RECT 72.225 91.075 72.395 91.245 ;
        RECT 72.685 91.075 72.855 91.245 ;
        RECT 73.145 91.075 73.315 91.245 ;
        RECT 73.605 91.075 73.775 91.245 ;
        RECT 74.065 91.075 74.235 91.245 ;
        RECT 74.525 91.075 74.695 91.245 ;
        RECT 74.985 91.075 75.155 91.245 ;
        RECT 75.445 91.075 75.615 91.245 ;
        RECT 75.905 91.075 76.075 91.245 ;
        RECT 76.365 91.075 76.535 91.245 ;
        RECT 76.825 91.075 76.995 91.245 ;
        RECT 77.285 91.075 77.455 91.245 ;
        RECT 77.745 91.075 77.915 91.245 ;
        RECT 78.205 91.075 78.375 91.245 ;
        RECT 78.665 91.075 78.835 91.245 ;
        RECT 79.125 91.075 79.295 91.245 ;
        RECT 79.585 91.075 79.755 91.245 ;
        RECT 80.045 91.075 80.215 91.245 ;
        RECT 80.505 91.075 80.675 91.245 ;
        RECT 80.965 91.075 81.135 91.245 ;
        RECT 81.425 91.075 81.595 91.245 ;
        RECT 81.885 91.075 82.055 91.245 ;
        RECT 82.345 91.075 82.515 91.245 ;
        RECT 82.805 91.075 82.975 91.245 ;
        RECT 83.265 91.075 83.435 91.245 ;
        RECT 83.725 91.075 83.895 91.245 ;
        RECT 84.185 91.075 84.355 91.245 ;
        RECT 84.645 91.075 84.815 91.245 ;
        RECT 85.105 91.075 85.275 91.245 ;
        RECT 85.565 91.075 85.735 91.245 ;
        RECT 86.025 91.075 86.195 91.245 ;
        RECT 86.485 91.075 86.655 91.245 ;
        RECT 86.945 91.075 87.115 91.245 ;
        RECT 87.405 91.075 87.575 91.245 ;
        RECT 87.865 91.075 88.035 91.245 ;
        RECT 88.325 91.075 88.495 91.245 ;
        RECT 88.785 91.075 88.955 91.245 ;
        RECT 89.245 91.075 89.415 91.245 ;
        RECT 89.705 91.075 89.875 91.245 ;
        RECT 90.165 91.075 90.335 91.245 ;
        RECT 90.625 91.075 90.795 91.245 ;
        RECT 91.085 91.075 91.255 91.245 ;
        RECT 91.545 91.075 91.715 91.245 ;
        RECT 92.005 91.075 92.175 91.245 ;
        RECT 92.465 91.075 92.635 91.245 ;
        RECT 92.925 91.075 93.095 91.245 ;
        RECT 93.385 91.075 93.555 91.245 ;
        RECT 93.845 91.075 94.015 91.245 ;
        RECT 94.305 91.075 94.475 91.245 ;
        RECT 94.765 91.075 94.935 91.245 ;
        RECT 95.225 91.075 95.395 91.245 ;
        RECT 95.685 91.075 95.855 91.245 ;
        RECT 96.145 91.075 96.315 91.245 ;
        RECT 96.605 91.075 96.775 91.245 ;
        RECT 97.065 91.075 97.235 91.245 ;
        RECT 97.525 91.075 97.695 91.245 ;
        RECT 97.985 91.075 98.155 91.245 ;
        RECT 98.445 91.075 98.615 91.245 ;
        RECT 98.905 91.075 99.075 91.245 ;
        RECT 99.365 91.075 99.535 91.245 ;
        RECT 99.825 91.075 99.995 91.245 ;
        RECT 100.285 91.075 100.455 91.245 ;
        RECT 100.745 91.075 100.915 91.245 ;
        RECT 101.205 91.075 101.375 91.245 ;
        RECT 101.665 91.075 101.835 91.245 ;
        RECT 102.125 91.075 102.295 91.245 ;
        RECT 102.585 91.075 102.755 91.245 ;
        RECT 103.045 91.075 103.215 91.245 ;
        RECT 103.505 91.075 103.675 91.245 ;
        RECT 103.965 91.075 104.135 91.245 ;
        RECT 104.425 91.075 104.595 91.245 ;
        RECT 104.885 91.075 105.055 91.245 ;
        RECT 105.345 91.075 105.515 91.245 ;
        RECT 105.805 91.075 105.975 91.245 ;
        RECT 106.265 91.075 106.435 91.245 ;
        RECT 106.725 91.075 106.895 91.245 ;
        RECT 107.185 91.075 107.355 91.245 ;
        RECT 107.645 91.075 107.815 91.245 ;
        RECT 108.105 91.075 108.275 91.245 ;
        RECT 108.565 91.075 108.735 91.245 ;
        RECT 109.025 91.075 109.195 91.245 ;
        RECT 109.485 91.075 109.655 91.245 ;
        RECT 109.945 91.075 110.115 91.245 ;
        RECT 110.405 91.075 110.575 91.245 ;
        RECT 110.865 91.075 111.035 91.245 ;
        RECT 111.325 91.075 111.495 91.245 ;
        RECT 111.785 91.075 111.955 91.245 ;
        RECT 112.245 91.075 112.415 91.245 ;
        RECT 112.705 91.075 112.875 91.245 ;
        RECT 113.165 91.075 113.335 91.245 ;
        RECT 113.625 91.075 113.795 91.245 ;
        RECT 114.085 91.075 114.255 91.245 ;
        RECT 114.545 91.075 114.715 91.245 ;
        RECT 115.005 91.075 115.175 91.245 ;
        RECT 115.465 91.075 115.635 91.245 ;
        RECT 115.925 91.075 116.095 91.245 ;
        RECT 116.385 91.075 116.555 91.245 ;
        RECT 116.845 91.075 117.015 91.245 ;
        RECT 117.305 91.075 117.475 91.245 ;
        RECT 117.765 91.075 117.935 91.245 ;
        RECT 118.225 91.075 118.395 91.245 ;
        RECT 118.685 91.075 118.855 91.245 ;
        RECT 119.145 91.075 119.315 91.245 ;
        RECT 119.605 91.075 119.775 91.245 ;
        RECT 120.065 91.075 120.235 91.245 ;
        RECT 120.525 91.075 120.695 91.245 ;
        RECT 120.985 91.075 121.155 91.245 ;
        RECT 121.445 91.075 121.615 91.245 ;
        RECT 121.905 91.075 122.075 91.245 ;
        RECT 122.365 91.075 122.535 91.245 ;
        RECT 122.825 91.075 122.995 91.245 ;
        RECT 123.285 91.075 123.455 91.245 ;
        RECT 123.745 91.075 123.915 91.245 ;
        RECT 124.205 91.075 124.375 91.245 ;
        RECT 124.665 91.075 124.835 91.245 ;
        RECT 125.125 91.075 125.295 91.245 ;
        RECT 125.585 91.075 125.755 91.245 ;
        RECT 126.045 91.075 126.215 91.245 ;
        RECT 126.505 91.075 126.675 91.245 ;
        RECT 126.965 91.075 127.135 91.245 ;
        RECT 127.425 91.075 127.595 91.245 ;
        RECT 127.885 91.075 128.055 91.245 ;
        RECT 128.345 91.075 128.515 91.245 ;
        RECT 128.805 91.075 128.975 91.245 ;
        RECT 129.265 91.075 129.435 91.245 ;
        RECT 129.725 91.075 129.895 91.245 ;
        RECT 130.185 91.075 130.355 91.245 ;
        RECT 130.645 91.075 130.815 91.245 ;
        RECT 131.105 91.075 131.275 91.245 ;
        RECT 131.565 91.075 131.735 91.245 ;
        RECT 132.025 91.075 132.195 91.245 ;
        RECT 132.485 91.075 132.655 91.245 ;
        RECT 132.945 91.075 133.115 91.245 ;
        RECT 133.405 91.075 133.575 91.245 ;
        RECT 133.865 91.075 134.035 91.245 ;
        RECT 134.325 91.075 134.495 91.245 ;
        RECT 134.785 91.075 134.955 91.245 ;
        RECT 135.245 91.075 135.415 91.245 ;
        RECT 135.705 91.075 135.875 91.245 ;
        RECT 136.165 91.075 136.335 91.245 ;
        RECT 136.625 91.075 136.795 91.245 ;
        RECT 137.085 91.075 137.255 91.245 ;
        RECT 137.545 91.075 137.715 91.245 ;
        RECT 138.005 91.075 138.175 91.245 ;
        RECT 138.465 91.075 138.635 91.245 ;
        RECT 138.925 91.075 139.095 91.245 ;
        RECT 139.385 91.075 139.555 91.245 ;
        RECT 139.845 91.075 140.015 91.245 ;
        RECT 140.305 91.075 140.475 91.245 ;
        RECT 140.765 91.075 140.935 91.245 ;
        RECT 141.225 91.075 141.395 91.245 ;
        RECT 141.685 91.075 141.855 91.245 ;
        RECT 142.145 91.075 142.315 91.245 ;
        RECT 142.605 91.075 142.775 91.245 ;
        RECT 143.065 91.075 143.235 91.245 ;
        RECT 143.525 91.075 143.695 91.245 ;
        RECT 143.985 91.075 144.155 91.245 ;
        RECT 55.665 85.635 55.835 85.805 ;
        RECT 56.125 85.635 56.295 85.805 ;
        RECT 56.585 85.635 56.755 85.805 ;
        RECT 57.045 85.635 57.215 85.805 ;
        RECT 57.505 85.635 57.675 85.805 ;
        RECT 57.965 85.635 58.135 85.805 ;
        RECT 58.425 85.635 58.595 85.805 ;
        RECT 58.885 85.635 59.055 85.805 ;
        RECT 59.345 85.635 59.515 85.805 ;
        RECT 59.805 85.635 59.975 85.805 ;
        RECT 60.265 85.635 60.435 85.805 ;
        RECT 60.725 85.635 60.895 85.805 ;
        RECT 61.185 85.635 61.355 85.805 ;
        RECT 61.645 85.635 61.815 85.805 ;
        RECT 62.105 85.635 62.275 85.805 ;
        RECT 62.565 85.635 62.735 85.805 ;
        RECT 63.025 85.635 63.195 85.805 ;
        RECT 63.485 85.635 63.655 85.805 ;
        RECT 63.945 85.635 64.115 85.805 ;
        RECT 64.405 85.635 64.575 85.805 ;
        RECT 64.865 85.635 65.035 85.805 ;
        RECT 65.325 85.635 65.495 85.805 ;
        RECT 65.785 85.635 65.955 85.805 ;
        RECT 66.245 85.635 66.415 85.805 ;
        RECT 66.705 85.635 66.875 85.805 ;
        RECT 67.165 85.635 67.335 85.805 ;
        RECT 67.625 85.635 67.795 85.805 ;
        RECT 68.085 85.635 68.255 85.805 ;
        RECT 68.545 85.635 68.715 85.805 ;
        RECT 69.005 85.635 69.175 85.805 ;
        RECT 69.465 85.635 69.635 85.805 ;
        RECT 69.925 85.635 70.095 85.805 ;
        RECT 70.385 85.635 70.555 85.805 ;
        RECT 70.845 85.635 71.015 85.805 ;
        RECT 71.305 85.635 71.475 85.805 ;
        RECT 71.765 85.635 71.935 85.805 ;
        RECT 72.225 85.635 72.395 85.805 ;
        RECT 72.685 85.635 72.855 85.805 ;
        RECT 73.145 85.635 73.315 85.805 ;
        RECT 73.605 85.635 73.775 85.805 ;
        RECT 74.065 85.635 74.235 85.805 ;
        RECT 74.525 85.635 74.695 85.805 ;
        RECT 74.985 85.635 75.155 85.805 ;
        RECT 75.445 85.635 75.615 85.805 ;
        RECT 75.905 85.635 76.075 85.805 ;
        RECT 76.365 85.635 76.535 85.805 ;
        RECT 76.825 85.635 76.995 85.805 ;
        RECT 77.285 85.635 77.455 85.805 ;
        RECT 77.745 85.635 77.915 85.805 ;
        RECT 78.205 85.635 78.375 85.805 ;
        RECT 78.665 85.635 78.835 85.805 ;
        RECT 79.125 85.635 79.295 85.805 ;
        RECT 79.585 85.635 79.755 85.805 ;
        RECT 80.045 85.635 80.215 85.805 ;
        RECT 80.505 85.635 80.675 85.805 ;
        RECT 80.965 85.635 81.135 85.805 ;
        RECT 81.425 85.635 81.595 85.805 ;
        RECT 81.885 85.635 82.055 85.805 ;
        RECT 82.345 85.635 82.515 85.805 ;
        RECT 82.805 85.635 82.975 85.805 ;
        RECT 83.265 85.635 83.435 85.805 ;
        RECT 83.725 85.635 83.895 85.805 ;
        RECT 84.185 85.635 84.355 85.805 ;
        RECT 84.645 85.635 84.815 85.805 ;
        RECT 85.105 85.635 85.275 85.805 ;
        RECT 85.565 85.635 85.735 85.805 ;
        RECT 86.025 85.635 86.195 85.805 ;
        RECT 86.485 85.635 86.655 85.805 ;
        RECT 86.945 85.635 87.115 85.805 ;
        RECT 87.405 85.635 87.575 85.805 ;
        RECT 87.865 85.635 88.035 85.805 ;
        RECT 88.325 85.635 88.495 85.805 ;
        RECT 88.785 85.635 88.955 85.805 ;
        RECT 89.245 85.635 89.415 85.805 ;
        RECT 89.705 85.635 89.875 85.805 ;
        RECT 90.165 85.635 90.335 85.805 ;
        RECT 90.625 85.635 90.795 85.805 ;
        RECT 91.085 85.635 91.255 85.805 ;
        RECT 91.545 85.635 91.715 85.805 ;
        RECT 92.005 85.635 92.175 85.805 ;
        RECT 92.465 85.635 92.635 85.805 ;
        RECT 92.925 85.635 93.095 85.805 ;
        RECT 93.385 85.635 93.555 85.805 ;
        RECT 93.845 85.635 94.015 85.805 ;
        RECT 94.305 85.635 94.475 85.805 ;
        RECT 94.765 85.635 94.935 85.805 ;
        RECT 95.225 85.635 95.395 85.805 ;
        RECT 95.685 85.635 95.855 85.805 ;
        RECT 96.145 85.635 96.315 85.805 ;
        RECT 96.605 85.635 96.775 85.805 ;
        RECT 97.065 85.635 97.235 85.805 ;
        RECT 97.525 85.635 97.695 85.805 ;
        RECT 97.985 85.635 98.155 85.805 ;
        RECT 98.445 85.635 98.615 85.805 ;
        RECT 98.905 85.635 99.075 85.805 ;
        RECT 99.365 85.635 99.535 85.805 ;
        RECT 99.825 85.635 99.995 85.805 ;
        RECT 100.285 85.635 100.455 85.805 ;
        RECT 100.745 85.635 100.915 85.805 ;
        RECT 101.205 85.635 101.375 85.805 ;
        RECT 101.665 85.635 101.835 85.805 ;
        RECT 102.125 85.635 102.295 85.805 ;
        RECT 102.585 85.635 102.755 85.805 ;
        RECT 103.045 85.635 103.215 85.805 ;
        RECT 103.505 85.635 103.675 85.805 ;
        RECT 103.965 85.635 104.135 85.805 ;
        RECT 104.425 85.635 104.595 85.805 ;
        RECT 104.885 85.635 105.055 85.805 ;
        RECT 105.345 85.635 105.515 85.805 ;
        RECT 105.805 85.635 105.975 85.805 ;
        RECT 106.265 85.635 106.435 85.805 ;
        RECT 106.725 85.635 106.895 85.805 ;
        RECT 107.185 85.635 107.355 85.805 ;
        RECT 107.645 85.635 107.815 85.805 ;
        RECT 108.105 85.635 108.275 85.805 ;
        RECT 108.565 85.635 108.735 85.805 ;
        RECT 109.025 85.635 109.195 85.805 ;
        RECT 109.485 85.635 109.655 85.805 ;
        RECT 109.945 85.635 110.115 85.805 ;
        RECT 110.405 85.635 110.575 85.805 ;
        RECT 110.865 85.635 111.035 85.805 ;
        RECT 111.325 85.635 111.495 85.805 ;
        RECT 111.785 85.635 111.955 85.805 ;
        RECT 112.245 85.635 112.415 85.805 ;
        RECT 112.705 85.635 112.875 85.805 ;
        RECT 113.165 85.635 113.335 85.805 ;
        RECT 113.625 85.635 113.795 85.805 ;
        RECT 114.085 85.635 114.255 85.805 ;
        RECT 114.545 85.635 114.715 85.805 ;
        RECT 115.005 85.635 115.175 85.805 ;
        RECT 115.465 85.635 115.635 85.805 ;
        RECT 115.925 85.635 116.095 85.805 ;
        RECT 116.385 85.635 116.555 85.805 ;
        RECT 116.845 85.635 117.015 85.805 ;
        RECT 117.305 85.635 117.475 85.805 ;
        RECT 117.765 85.635 117.935 85.805 ;
        RECT 118.225 85.635 118.395 85.805 ;
        RECT 118.685 85.635 118.855 85.805 ;
        RECT 119.145 85.635 119.315 85.805 ;
        RECT 119.605 85.635 119.775 85.805 ;
        RECT 120.065 85.635 120.235 85.805 ;
        RECT 120.525 85.635 120.695 85.805 ;
        RECT 120.985 85.635 121.155 85.805 ;
        RECT 121.445 85.635 121.615 85.805 ;
        RECT 121.905 85.635 122.075 85.805 ;
        RECT 122.365 85.635 122.535 85.805 ;
        RECT 122.825 85.635 122.995 85.805 ;
        RECT 123.285 85.635 123.455 85.805 ;
        RECT 123.745 85.635 123.915 85.805 ;
        RECT 124.205 85.635 124.375 85.805 ;
        RECT 124.665 85.635 124.835 85.805 ;
        RECT 125.125 85.635 125.295 85.805 ;
        RECT 125.585 85.635 125.755 85.805 ;
        RECT 126.045 85.635 126.215 85.805 ;
        RECT 126.505 85.635 126.675 85.805 ;
        RECT 126.965 85.635 127.135 85.805 ;
        RECT 127.425 85.635 127.595 85.805 ;
        RECT 127.885 85.635 128.055 85.805 ;
        RECT 128.345 85.635 128.515 85.805 ;
        RECT 128.805 85.635 128.975 85.805 ;
        RECT 129.265 85.635 129.435 85.805 ;
        RECT 129.725 85.635 129.895 85.805 ;
        RECT 130.185 85.635 130.355 85.805 ;
        RECT 130.645 85.635 130.815 85.805 ;
        RECT 131.105 85.635 131.275 85.805 ;
        RECT 131.565 85.635 131.735 85.805 ;
        RECT 132.025 85.635 132.195 85.805 ;
        RECT 132.485 85.635 132.655 85.805 ;
        RECT 132.945 85.635 133.115 85.805 ;
        RECT 133.405 85.635 133.575 85.805 ;
        RECT 133.865 85.635 134.035 85.805 ;
        RECT 134.325 85.635 134.495 85.805 ;
        RECT 134.785 85.635 134.955 85.805 ;
        RECT 135.245 85.635 135.415 85.805 ;
        RECT 135.705 85.635 135.875 85.805 ;
        RECT 136.165 85.635 136.335 85.805 ;
        RECT 136.625 85.635 136.795 85.805 ;
        RECT 137.085 85.635 137.255 85.805 ;
        RECT 137.545 85.635 137.715 85.805 ;
        RECT 138.005 85.635 138.175 85.805 ;
        RECT 138.465 85.635 138.635 85.805 ;
        RECT 138.925 85.635 139.095 85.805 ;
        RECT 139.385 85.635 139.555 85.805 ;
        RECT 139.845 85.635 140.015 85.805 ;
        RECT 140.305 85.635 140.475 85.805 ;
        RECT 140.765 85.635 140.935 85.805 ;
        RECT 141.225 85.635 141.395 85.805 ;
        RECT 141.685 85.635 141.855 85.805 ;
        RECT 142.145 85.635 142.315 85.805 ;
        RECT 142.605 85.635 142.775 85.805 ;
        RECT 143.065 85.635 143.235 85.805 ;
        RECT 143.525 85.635 143.695 85.805 ;
        RECT 143.985 85.635 144.155 85.805 ;
        RECT 55.665 80.195 55.835 80.365 ;
        RECT 56.125 80.195 56.295 80.365 ;
        RECT 56.585 80.195 56.755 80.365 ;
        RECT 57.045 80.195 57.215 80.365 ;
        RECT 57.505 80.195 57.675 80.365 ;
        RECT 57.965 80.195 58.135 80.365 ;
        RECT 58.425 80.195 58.595 80.365 ;
        RECT 58.885 80.195 59.055 80.365 ;
        RECT 59.345 80.195 59.515 80.365 ;
        RECT 59.805 80.195 59.975 80.365 ;
        RECT 60.265 80.195 60.435 80.365 ;
        RECT 60.725 80.195 60.895 80.365 ;
        RECT 61.185 80.195 61.355 80.365 ;
        RECT 61.645 80.195 61.815 80.365 ;
        RECT 62.105 80.195 62.275 80.365 ;
        RECT 62.565 80.195 62.735 80.365 ;
        RECT 63.025 80.195 63.195 80.365 ;
        RECT 63.485 80.195 63.655 80.365 ;
        RECT 63.945 80.195 64.115 80.365 ;
        RECT 64.405 80.195 64.575 80.365 ;
        RECT 64.865 80.195 65.035 80.365 ;
        RECT 65.325 80.195 65.495 80.365 ;
        RECT 65.785 80.195 65.955 80.365 ;
        RECT 66.245 80.195 66.415 80.365 ;
        RECT 66.705 80.195 66.875 80.365 ;
        RECT 67.165 80.195 67.335 80.365 ;
        RECT 67.625 80.195 67.795 80.365 ;
        RECT 68.085 80.195 68.255 80.365 ;
        RECT 68.545 80.195 68.715 80.365 ;
        RECT 69.005 80.195 69.175 80.365 ;
        RECT 69.465 80.195 69.635 80.365 ;
        RECT 69.925 80.195 70.095 80.365 ;
        RECT 70.385 80.195 70.555 80.365 ;
        RECT 70.845 80.195 71.015 80.365 ;
        RECT 71.305 80.195 71.475 80.365 ;
        RECT 71.765 80.195 71.935 80.365 ;
        RECT 72.225 80.195 72.395 80.365 ;
        RECT 72.685 80.195 72.855 80.365 ;
        RECT 73.145 80.195 73.315 80.365 ;
        RECT 73.605 80.195 73.775 80.365 ;
        RECT 74.065 80.195 74.235 80.365 ;
        RECT 74.525 80.195 74.695 80.365 ;
        RECT 74.985 80.195 75.155 80.365 ;
        RECT 75.445 80.195 75.615 80.365 ;
        RECT 75.905 80.195 76.075 80.365 ;
        RECT 76.365 80.195 76.535 80.365 ;
        RECT 76.825 80.195 76.995 80.365 ;
        RECT 77.285 80.195 77.455 80.365 ;
        RECT 77.745 80.195 77.915 80.365 ;
        RECT 78.205 80.195 78.375 80.365 ;
        RECT 78.665 80.195 78.835 80.365 ;
        RECT 79.125 80.195 79.295 80.365 ;
        RECT 79.585 80.195 79.755 80.365 ;
        RECT 80.045 80.195 80.215 80.365 ;
        RECT 80.505 80.195 80.675 80.365 ;
        RECT 80.965 80.195 81.135 80.365 ;
        RECT 81.425 80.195 81.595 80.365 ;
        RECT 81.885 80.195 82.055 80.365 ;
        RECT 82.345 80.195 82.515 80.365 ;
        RECT 82.805 80.195 82.975 80.365 ;
        RECT 83.265 80.195 83.435 80.365 ;
        RECT 83.725 80.195 83.895 80.365 ;
        RECT 84.185 80.195 84.355 80.365 ;
        RECT 84.645 80.195 84.815 80.365 ;
        RECT 85.105 80.195 85.275 80.365 ;
        RECT 85.565 80.195 85.735 80.365 ;
        RECT 86.025 80.195 86.195 80.365 ;
        RECT 86.485 80.195 86.655 80.365 ;
        RECT 86.945 80.195 87.115 80.365 ;
        RECT 87.405 80.195 87.575 80.365 ;
        RECT 87.865 80.195 88.035 80.365 ;
        RECT 88.325 80.195 88.495 80.365 ;
        RECT 88.785 80.195 88.955 80.365 ;
        RECT 89.245 80.195 89.415 80.365 ;
        RECT 89.705 80.195 89.875 80.365 ;
        RECT 90.165 80.195 90.335 80.365 ;
        RECT 90.625 80.195 90.795 80.365 ;
        RECT 91.085 80.195 91.255 80.365 ;
        RECT 91.545 80.195 91.715 80.365 ;
        RECT 92.005 80.195 92.175 80.365 ;
        RECT 92.465 80.195 92.635 80.365 ;
        RECT 92.925 80.195 93.095 80.365 ;
        RECT 93.385 80.195 93.555 80.365 ;
        RECT 93.845 80.195 94.015 80.365 ;
        RECT 94.305 80.195 94.475 80.365 ;
        RECT 94.765 80.195 94.935 80.365 ;
        RECT 95.225 80.195 95.395 80.365 ;
        RECT 95.685 80.195 95.855 80.365 ;
        RECT 96.145 80.195 96.315 80.365 ;
        RECT 96.605 80.195 96.775 80.365 ;
        RECT 97.065 80.195 97.235 80.365 ;
        RECT 97.525 80.195 97.695 80.365 ;
        RECT 97.985 80.195 98.155 80.365 ;
        RECT 98.445 80.195 98.615 80.365 ;
        RECT 98.905 80.195 99.075 80.365 ;
        RECT 99.365 80.195 99.535 80.365 ;
        RECT 99.825 80.195 99.995 80.365 ;
        RECT 100.285 80.195 100.455 80.365 ;
        RECT 100.745 80.195 100.915 80.365 ;
        RECT 101.205 80.195 101.375 80.365 ;
        RECT 101.665 80.195 101.835 80.365 ;
        RECT 102.125 80.195 102.295 80.365 ;
        RECT 102.585 80.195 102.755 80.365 ;
        RECT 103.045 80.195 103.215 80.365 ;
        RECT 103.505 80.195 103.675 80.365 ;
        RECT 103.965 80.195 104.135 80.365 ;
        RECT 104.425 80.195 104.595 80.365 ;
        RECT 104.885 80.195 105.055 80.365 ;
        RECT 105.345 80.195 105.515 80.365 ;
        RECT 105.805 80.195 105.975 80.365 ;
        RECT 106.265 80.195 106.435 80.365 ;
        RECT 106.725 80.195 106.895 80.365 ;
        RECT 107.185 80.195 107.355 80.365 ;
        RECT 107.645 80.195 107.815 80.365 ;
        RECT 108.105 80.195 108.275 80.365 ;
        RECT 108.565 80.195 108.735 80.365 ;
        RECT 109.025 80.195 109.195 80.365 ;
        RECT 109.485 80.195 109.655 80.365 ;
        RECT 109.945 80.195 110.115 80.365 ;
        RECT 110.405 80.195 110.575 80.365 ;
        RECT 110.865 80.195 111.035 80.365 ;
        RECT 111.325 80.195 111.495 80.365 ;
        RECT 111.785 80.195 111.955 80.365 ;
        RECT 112.245 80.195 112.415 80.365 ;
        RECT 112.705 80.195 112.875 80.365 ;
        RECT 113.165 80.195 113.335 80.365 ;
        RECT 113.625 80.195 113.795 80.365 ;
        RECT 114.085 80.195 114.255 80.365 ;
        RECT 114.545 80.195 114.715 80.365 ;
        RECT 115.005 80.195 115.175 80.365 ;
        RECT 115.465 80.195 115.635 80.365 ;
        RECT 115.925 80.195 116.095 80.365 ;
        RECT 116.385 80.195 116.555 80.365 ;
        RECT 116.845 80.195 117.015 80.365 ;
        RECT 117.305 80.195 117.475 80.365 ;
        RECT 117.765 80.195 117.935 80.365 ;
        RECT 118.225 80.195 118.395 80.365 ;
        RECT 118.685 80.195 118.855 80.365 ;
        RECT 119.145 80.195 119.315 80.365 ;
        RECT 119.605 80.195 119.775 80.365 ;
        RECT 120.065 80.195 120.235 80.365 ;
        RECT 120.525 80.195 120.695 80.365 ;
        RECT 120.985 80.195 121.155 80.365 ;
        RECT 121.445 80.195 121.615 80.365 ;
        RECT 121.905 80.195 122.075 80.365 ;
        RECT 122.365 80.195 122.535 80.365 ;
        RECT 122.825 80.195 122.995 80.365 ;
        RECT 123.285 80.195 123.455 80.365 ;
        RECT 123.745 80.195 123.915 80.365 ;
        RECT 124.205 80.195 124.375 80.365 ;
        RECT 124.665 80.195 124.835 80.365 ;
        RECT 125.125 80.195 125.295 80.365 ;
        RECT 125.585 80.195 125.755 80.365 ;
        RECT 126.045 80.195 126.215 80.365 ;
        RECT 126.505 80.195 126.675 80.365 ;
        RECT 126.965 80.195 127.135 80.365 ;
        RECT 127.425 80.195 127.595 80.365 ;
        RECT 127.885 80.195 128.055 80.365 ;
        RECT 128.345 80.195 128.515 80.365 ;
        RECT 128.805 80.195 128.975 80.365 ;
        RECT 129.265 80.195 129.435 80.365 ;
        RECT 129.725 80.195 129.895 80.365 ;
        RECT 130.185 80.195 130.355 80.365 ;
        RECT 130.645 80.195 130.815 80.365 ;
        RECT 131.105 80.195 131.275 80.365 ;
        RECT 131.565 80.195 131.735 80.365 ;
        RECT 132.025 80.195 132.195 80.365 ;
        RECT 132.485 80.195 132.655 80.365 ;
        RECT 132.945 80.195 133.115 80.365 ;
        RECT 133.405 80.195 133.575 80.365 ;
        RECT 133.865 80.195 134.035 80.365 ;
        RECT 134.325 80.195 134.495 80.365 ;
        RECT 134.785 80.195 134.955 80.365 ;
        RECT 135.245 80.195 135.415 80.365 ;
        RECT 135.705 80.195 135.875 80.365 ;
        RECT 136.165 80.195 136.335 80.365 ;
        RECT 136.625 80.195 136.795 80.365 ;
        RECT 137.085 80.195 137.255 80.365 ;
        RECT 137.545 80.195 137.715 80.365 ;
        RECT 138.005 80.195 138.175 80.365 ;
        RECT 138.465 80.195 138.635 80.365 ;
        RECT 138.925 80.195 139.095 80.365 ;
        RECT 139.385 80.195 139.555 80.365 ;
        RECT 139.845 80.195 140.015 80.365 ;
        RECT 140.305 80.195 140.475 80.365 ;
        RECT 140.765 80.195 140.935 80.365 ;
        RECT 141.225 80.195 141.395 80.365 ;
        RECT 141.685 80.195 141.855 80.365 ;
        RECT 142.145 80.195 142.315 80.365 ;
        RECT 142.605 80.195 142.775 80.365 ;
        RECT 143.065 80.195 143.235 80.365 ;
        RECT 143.525 80.195 143.695 80.365 ;
        RECT 143.985 80.195 144.155 80.365 ;
        RECT 55.665 74.755 55.835 74.925 ;
        RECT 56.125 74.755 56.295 74.925 ;
        RECT 56.585 74.755 56.755 74.925 ;
        RECT 57.045 74.755 57.215 74.925 ;
        RECT 57.505 74.755 57.675 74.925 ;
        RECT 57.965 74.755 58.135 74.925 ;
        RECT 58.425 74.755 58.595 74.925 ;
        RECT 58.885 74.755 59.055 74.925 ;
        RECT 59.345 74.755 59.515 74.925 ;
        RECT 59.805 74.755 59.975 74.925 ;
        RECT 60.265 74.755 60.435 74.925 ;
        RECT 60.725 74.755 60.895 74.925 ;
        RECT 61.185 74.755 61.355 74.925 ;
        RECT 61.645 74.755 61.815 74.925 ;
        RECT 62.105 74.755 62.275 74.925 ;
        RECT 62.565 74.755 62.735 74.925 ;
        RECT 63.025 74.755 63.195 74.925 ;
        RECT 63.485 74.755 63.655 74.925 ;
        RECT 63.945 74.755 64.115 74.925 ;
        RECT 64.405 74.755 64.575 74.925 ;
        RECT 64.865 74.755 65.035 74.925 ;
        RECT 65.325 74.755 65.495 74.925 ;
        RECT 65.785 74.755 65.955 74.925 ;
        RECT 66.245 74.755 66.415 74.925 ;
        RECT 66.705 74.755 66.875 74.925 ;
        RECT 67.165 74.755 67.335 74.925 ;
        RECT 67.625 74.755 67.795 74.925 ;
        RECT 68.085 74.755 68.255 74.925 ;
        RECT 68.545 74.755 68.715 74.925 ;
        RECT 69.005 74.755 69.175 74.925 ;
        RECT 69.465 74.755 69.635 74.925 ;
        RECT 69.925 74.755 70.095 74.925 ;
        RECT 70.385 74.755 70.555 74.925 ;
        RECT 70.845 74.755 71.015 74.925 ;
        RECT 71.305 74.755 71.475 74.925 ;
        RECT 71.765 74.755 71.935 74.925 ;
        RECT 72.225 74.755 72.395 74.925 ;
        RECT 72.685 74.755 72.855 74.925 ;
        RECT 73.145 74.755 73.315 74.925 ;
        RECT 73.605 74.755 73.775 74.925 ;
        RECT 74.065 74.755 74.235 74.925 ;
        RECT 74.525 74.755 74.695 74.925 ;
        RECT 74.985 74.755 75.155 74.925 ;
        RECT 75.445 74.755 75.615 74.925 ;
        RECT 75.905 74.755 76.075 74.925 ;
        RECT 76.365 74.755 76.535 74.925 ;
        RECT 76.825 74.755 76.995 74.925 ;
        RECT 77.285 74.755 77.455 74.925 ;
        RECT 77.745 74.755 77.915 74.925 ;
        RECT 78.205 74.755 78.375 74.925 ;
        RECT 78.665 74.755 78.835 74.925 ;
        RECT 79.125 74.755 79.295 74.925 ;
        RECT 79.585 74.755 79.755 74.925 ;
        RECT 80.045 74.755 80.215 74.925 ;
        RECT 80.505 74.755 80.675 74.925 ;
        RECT 80.965 74.755 81.135 74.925 ;
        RECT 81.425 74.755 81.595 74.925 ;
        RECT 81.885 74.755 82.055 74.925 ;
        RECT 82.345 74.755 82.515 74.925 ;
        RECT 82.805 74.755 82.975 74.925 ;
        RECT 83.265 74.755 83.435 74.925 ;
        RECT 83.725 74.755 83.895 74.925 ;
        RECT 84.185 74.755 84.355 74.925 ;
        RECT 84.645 74.755 84.815 74.925 ;
        RECT 85.105 74.755 85.275 74.925 ;
        RECT 85.565 74.755 85.735 74.925 ;
        RECT 86.025 74.755 86.195 74.925 ;
        RECT 86.485 74.755 86.655 74.925 ;
        RECT 86.945 74.755 87.115 74.925 ;
        RECT 87.405 74.755 87.575 74.925 ;
        RECT 87.865 74.755 88.035 74.925 ;
        RECT 88.325 74.755 88.495 74.925 ;
        RECT 88.785 74.755 88.955 74.925 ;
        RECT 89.245 74.755 89.415 74.925 ;
        RECT 89.705 74.755 89.875 74.925 ;
        RECT 90.165 74.755 90.335 74.925 ;
        RECT 90.625 74.755 90.795 74.925 ;
        RECT 91.085 74.755 91.255 74.925 ;
        RECT 91.545 74.755 91.715 74.925 ;
        RECT 92.005 74.755 92.175 74.925 ;
        RECT 92.465 74.755 92.635 74.925 ;
        RECT 92.925 74.755 93.095 74.925 ;
        RECT 93.385 74.755 93.555 74.925 ;
        RECT 93.845 74.755 94.015 74.925 ;
        RECT 94.305 74.755 94.475 74.925 ;
        RECT 94.765 74.755 94.935 74.925 ;
        RECT 95.225 74.755 95.395 74.925 ;
        RECT 95.685 74.755 95.855 74.925 ;
        RECT 96.145 74.755 96.315 74.925 ;
        RECT 96.605 74.755 96.775 74.925 ;
        RECT 97.065 74.755 97.235 74.925 ;
        RECT 97.525 74.755 97.695 74.925 ;
        RECT 97.985 74.755 98.155 74.925 ;
        RECT 98.445 74.755 98.615 74.925 ;
        RECT 98.905 74.755 99.075 74.925 ;
        RECT 99.365 74.755 99.535 74.925 ;
        RECT 99.825 74.755 99.995 74.925 ;
        RECT 100.285 74.755 100.455 74.925 ;
        RECT 100.745 74.755 100.915 74.925 ;
        RECT 101.205 74.755 101.375 74.925 ;
        RECT 101.665 74.755 101.835 74.925 ;
        RECT 102.125 74.755 102.295 74.925 ;
        RECT 102.585 74.755 102.755 74.925 ;
        RECT 103.045 74.755 103.215 74.925 ;
        RECT 103.505 74.755 103.675 74.925 ;
        RECT 103.965 74.755 104.135 74.925 ;
        RECT 104.425 74.755 104.595 74.925 ;
        RECT 104.885 74.755 105.055 74.925 ;
        RECT 105.345 74.755 105.515 74.925 ;
        RECT 105.805 74.755 105.975 74.925 ;
        RECT 106.265 74.755 106.435 74.925 ;
        RECT 106.725 74.755 106.895 74.925 ;
        RECT 107.185 74.755 107.355 74.925 ;
        RECT 107.645 74.755 107.815 74.925 ;
        RECT 108.105 74.755 108.275 74.925 ;
        RECT 108.565 74.755 108.735 74.925 ;
        RECT 109.025 74.755 109.195 74.925 ;
        RECT 109.485 74.755 109.655 74.925 ;
        RECT 109.945 74.755 110.115 74.925 ;
        RECT 110.405 74.755 110.575 74.925 ;
        RECT 110.865 74.755 111.035 74.925 ;
        RECT 111.325 74.755 111.495 74.925 ;
        RECT 111.785 74.755 111.955 74.925 ;
        RECT 112.245 74.755 112.415 74.925 ;
        RECT 112.705 74.755 112.875 74.925 ;
        RECT 113.165 74.755 113.335 74.925 ;
        RECT 113.625 74.755 113.795 74.925 ;
        RECT 114.085 74.755 114.255 74.925 ;
        RECT 114.545 74.755 114.715 74.925 ;
        RECT 115.005 74.755 115.175 74.925 ;
        RECT 115.465 74.755 115.635 74.925 ;
        RECT 115.925 74.755 116.095 74.925 ;
        RECT 116.385 74.755 116.555 74.925 ;
        RECT 116.845 74.755 117.015 74.925 ;
        RECT 117.305 74.755 117.475 74.925 ;
        RECT 117.765 74.755 117.935 74.925 ;
        RECT 118.225 74.755 118.395 74.925 ;
        RECT 118.685 74.755 118.855 74.925 ;
        RECT 119.145 74.755 119.315 74.925 ;
        RECT 119.605 74.755 119.775 74.925 ;
        RECT 120.065 74.755 120.235 74.925 ;
        RECT 120.525 74.755 120.695 74.925 ;
        RECT 120.985 74.755 121.155 74.925 ;
        RECT 121.445 74.755 121.615 74.925 ;
        RECT 121.905 74.755 122.075 74.925 ;
        RECT 122.365 74.755 122.535 74.925 ;
        RECT 122.825 74.755 122.995 74.925 ;
        RECT 123.285 74.755 123.455 74.925 ;
        RECT 123.745 74.755 123.915 74.925 ;
        RECT 124.205 74.755 124.375 74.925 ;
        RECT 124.665 74.755 124.835 74.925 ;
        RECT 125.125 74.755 125.295 74.925 ;
        RECT 125.585 74.755 125.755 74.925 ;
        RECT 126.045 74.755 126.215 74.925 ;
        RECT 126.505 74.755 126.675 74.925 ;
        RECT 126.965 74.755 127.135 74.925 ;
        RECT 127.425 74.755 127.595 74.925 ;
        RECT 127.885 74.755 128.055 74.925 ;
        RECT 128.345 74.755 128.515 74.925 ;
        RECT 128.805 74.755 128.975 74.925 ;
        RECT 129.265 74.755 129.435 74.925 ;
        RECT 129.725 74.755 129.895 74.925 ;
        RECT 130.185 74.755 130.355 74.925 ;
        RECT 130.645 74.755 130.815 74.925 ;
        RECT 131.105 74.755 131.275 74.925 ;
        RECT 131.565 74.755 131.735 74.925 ;
        RECT 132.025 74.755 132.195 74.925 ;
        RECT 132.485 74.755 132.655 74.925 ;
        RECT 132.945 74.755 133.115 74.925 ;
        RECT 133.405 74.755 133.575 74.925 ;
        RECT 133.865 74.755 134.035 74.925 ;
        RECT 134.325 74.755 134.495 74.925 ;
        RECT 134.785 74.755 134.955 74.925 ;
        RECT 135.245 74.755 135.415 74.925 ;
        RECT 135.705 74.755 135.875 74.925 ;
        RECT 136.165 74.755 136.335 74.925 ;
        RECT 136.625 74.755 136.795 74.925 ;
        RECT 137.085 74.755 137.255 74.925 ;
        RECT 137.545 74.755 137.715 74.925 ;
        RECT 138.005 74.755 138.175 74.925 ;
        RECT 138.465 74.755 138.635 74.925 ;
        RECT 138.925 74.755 139.095 74.925 ;
        RECT 139.385 74.755 139.555 74.925 ;
        RECT 139.845 74.755 140.015 74.925 ;
        RECT 140.305 74.755 140.475 74.925 ;
        RECT 140.765 74.755 140.935 74.925 ;
        RECT 141.225 74.755 141.395 74.925 ;
        RECT 141.685 74.755 141.855 74.925 ;
        RECT 142.145 74.755 142.315 74.925 ;
        RECT 142.605 74.755 142.775 74.925 ;
        RECT 143.065 74.755 143.235 74.925 ;
        RECT 143.525 74.755 143.695 74.925 ;
        RECT 143.985 74.755 144.155 74.925 ;
        RECT 55.665 69.315 55.835 69.485 ;
        RECT 56.125 69.315 56.295 69.485 ;
        RECT 56.585 69.315 56.755 69.485 ;
        RECT 57.045 69.315 57.215 69.485 ;
        RECT 57.505 69.315 57.675 69.485 ;
        RECT 57.965 69.315 58.135 69.485 ;
        RECT 58.425 69.315 58.595 69.485 ;
        RECT 58.885 69.315 59.055 69.485 ;
        RECT 59.345 69.315 59.515 69.485 ;
        RECT 59.805 69.315 59.975 69.485 ;
        RECT 60.265 69.315 60.435 69.485 ;
        RECT 60.725 69.315 60.895 69.485 ;
        RECT 61.185 69.315 61.355 69.485 ;
        RECT 61.645 69.315 61.815 69.485 ;
        RECT 62.105 69.315 62.275 69.485 ;
        RECT 62.565 69.315 62.735 69.485 ;
        RECT 63.025 69.315 63.195 69.485 ;
        RECT 63.485 69.315 63.655 69.485 ;
        RECT 63.945 69.315 64.115 69.485 ;
        RECT 64.405 69.315 64.575 69.485 ;
        RECT 64.865 69.315 65.035 69.485 ;
        RECT 65.325 69.315 65.495 69.485 ;
        RECT 65.785 69.315 65.955 69.485 ;
        RECT 66.245 69.315 66.415 69.485 ;
        RECT 66.705 69.315 66.875 69.485 ;
        RECT 67.165 69.315 67.335 69.485 ;
        RECT 67.625 69.315 67.795 69.485 ;
        RECT 68.085 69.315 68.255 69.485 ;
        RECT 68.545 69.315 68.715 69.485 ;
        RECT 69.005 69.315 69.175 69.485 ;
        RECT 69.465 69.315 69.635 69.485 ;
        RECT 69.925 69.315 70.095 69.485 ;
        RECT 70.385 69.315 70.555 69.485 ;
        RECT 70.845 69.315 71.015 69.485 ;
        RECT 71.305 69.315 71.475 69.485 ;
        RECT 71.765 69.315 71.935 69.485 ;
        RECT 72.225 69.315 72.395 69.485 ;
        RECT 72.685 69.315 72.855 69.485 ;
        RECT 73.145 69.315 73.315 69.485 ;
        RECT 73.605 69.315 73.775 69.485 ;
        RECT 74.065 69.315 74.235 69.485 ;
        RECT 74.525 69.315 74.695 69.485 ;
        RECT 74.985 69.315 75.155 69.485 ;
        RECT 75.445 69.315 75.615 69.485 ;
        RECT 75.905 69.315 76.075 69.485 ;
        RECT 76.365 69.315 76.535 69.485 ;
        RECT 76.825 69.315 76.995 69.485 ;
        RECT 77.285 69.315 77.455 69.485 ;
        RECT 77.745 69.315 77.915 69.485 ;
        RECT 78.205 69.315 78.375 69.485 ;
        RECT 78.665 69.315 78.835 69.485 ;
        RECT 79.125 69.315 79.295 69.485 ;
        RECT 79.585 69.315 79.755 69.485 ;
        RECT 80.045 69.315 80.215 69.485 ;
        RECT 80.505 69.315 80.675 69.485 ;
        RECT 80.965 69.315 81.135 69.485 ;
        RECT 81.425 69.315 81.595 69.485 ;
        RECT 81.885 69.315 82.055 69.485 ;
        RECT 82.345 69.315 82.515 69.485 ;
        RECT 82.805 69.315 82.975 69.485 ;
        RECT 83.265 69.315 83.435 69.485 ;
        RECT 83.725 69.315 83.895 69.485 ;
        RECT 84.185 69.315 84.355 69.485 ;
        RECT 84.645 69.315 84.815 69.485 ;
        RECT 85.105 69.315 85.275 69.485 ;
        RECT 85.565 69.315 85.735 69.485 ;
        RECT 86.025 69.315 86.195 69.485 ;
        RECT 86.485 69.315 86.655 69.485 ;
        RECT 86.945 69.315 87.115 69.485 ;
        RECT 87.405 69.315 87.575 69.485 ;
        RECT 87.865 69.315 88.035 69.485 ;
        RECT 88.325 69.315 88.495 69.485 ;
        RECT 88.785 69.315 88.955 69.485 ;
        RECT 89.245 69.315 89.415 69.485 ;
        RECT 89.705 69.315 89.875 69.485 ;
        RECT 90.165 69.315 90.335 69.485 ;
        RECT 90.625 69.315 90.795 69.485 ;
        RECT 91.085 69.315 91.255 69.485 ;
        RECT 91.545 69.315 91.715 69.485 ;
        RECT 92.005 69.315 92.175 69.485 ;
        RECT 92.465 69.315 92.635 69.485 ;
        RECT 92.925 69.315 93.095 69.485 ;
        RECT 93.385 69.315 93.555 69.485 ;
        RECT 93.845 69.315 94.015 69.485 ;
        RECT 94.305 69.315 94.475 69.485 ;
        RECT 94.765 69.315 94.935 69.485 ;
        RECT 95.225 69.315 95.395 69.485 ;
        RECT 95.685 69.315 95.855 69.485 ;
        RECT 96.145 69.315 96.315 69.485 ;
        RECT 96.605 69.315 96.775 69.485 ;
        RECT 97.065 69.315 97.235 69.485 ;
        RECT 97.525 69.315 97.695 69.485 ;
        RECT 97.985 69.315 98.155 69.485 ;
        RECT 98.445 69.315 98.615 69.485 ;
        RECT 98.905 69.315 99.075 69.485 ;
        RECT 99.365 69.315 99.535 69.485 ;
        RECT 99.825 69.315 99.995 69.485 ;
        RECT 100.285 69.315 100.455 69.485 ;
        RECT 100.745 69.315 100.915 69.485 ;
        RECT 101.205 69.315 101.375 69.485 ;
        RECT 101.665 69.315 101.835 69.485 ;
        RECT 102.125 69.315 102.295 69.485 ;
        RECT 102.585 69.315 102.755 69.485 ;
        RECT 103.045 69.315 103.215 69.485 ;
        RECT 103.505 69.315 103.675 69.485 ;
        RECT 103.965 69.315 104.135 69.485 ;
        RECT 104.425 69.315 104.595 69.485 ;
        RECT 104.885 69.315 105.055 69.485 ;
        RECT 105.345 69.315 105.515 69.485 ;
        RECT 105.805 69.315 105.975 69.485 ;
        RECT 106.265 69.315 106.435 69.485 ;
        RECT 106.725 69.315 106.895 69.485 ;
        RECT 107.185 69.315 107.355 69.485 ;
        RECT 107.645 69.315 107.815 69.485 ;
        RECT 108.105 69.315 108.275 69.485 ;
        RECT 108.565 69.315 108.735 69.485 ;
        RECT 109.025 69.315 109.195 69.485 ;
        RECT 109.485 69.315 109.655 69.485 ;
        RECT 109.945 69.315 110.115 69.485 ;
        RECT 110.405 69.315 110.575 69.485 ;
        RECT 110.865 69.315 111.035 69.485 ;
        RECT 111.325 69.315 111.495 69.485 ;
        RECT 111.785 69.315 111.955 69.485 ;
        RECT 112.245 69.315 112.415 69.485 ;
        RECT 112.705 69.315 112.875 69.485 ;
        RECT 113.165 69.315 113.335 69.485 ;
        RECT 113.625 69.315 113.795 69.485 ;
        RECT 114.085 69.315 114.255 69.485 ;
        RECT 114.545 69.315 114.715 69.485 ;
        RECT 115.005 69.315 115.175 69.485 ;
        RECT 115.465 69.315 115.635 69.485 ;
        RECT 115.925 69.315 116.095 69.485 ;
        RECT 116.385 69.315 116.555 69.485 ;
        RECT 116.845 69.315 117.015 69.485 ;
        RECT 117.305 69.315 117.475 69.485 ;
        RECT 117.765 69.315 117.935 69.485 ;
        RECT 118.225 69.315 118.395 69.485 ;
        RECT 118.685 69.315 118.855 69.485 ;
        RECT 119.145 69.315 119.315 69.485 ;
        RECT 119.605 69.315 119.775 69.485 ;
        RECT 120.065 69.315 120.235 69.485 ;
        RECT 120.525 69.315 120.695 69.485 ;
        RECT 120.985 69.315 121.155 69.485 ;
        RECT 121.445 69.315 121.615 69.485 ;
        RECT 121.905 69.315 122.075 69.485 ;
        RECT 122.365 69.315 122.535 69.485 ;
        RECT 122.825 69.315 122.995 69.485 ;
        RECT 123.285 69.315 123.455 69.485 ;
        RECT 123.745 69.315 123.915 69.485 ;
        RECT 124.205 69.315 124.375 69.485 ;
        RECT 124.665 69.315 124.835 69.485 ;
        RECT 125.125 69.315 125.295 69.485 ;
        RECT 125.585 69.315 125.755 69.485 ;
        RECT 126.045 69.315 126.215 69.485 ;
        RECT 126.505 69.315 126.675 69.485 ;
        RECT 126.965 69.315 127.135 69.485 ;
        RECT 127.425 69.315 127.595 69.485 ;
        RECT 127.885 69.315 128.055 69.485 ;
        RECT 128.345 69.315 128.515 69.485 ;
        RECT 128.805 69.315 128.975 69.485 ;
        RECT 129.265 69.315 129.435 69.485 ;
        RECT 129.725 69.315 129.895 69.485 ;
        RECT 130.185 69.315 130.355 69.485 ;
        RECT 130.645 69.315 130.815 69.485 ;
        RECT 131.105 69.315 131.275 69.485 ;
        RECT 131.565 69.315 131.735 69.485 ;
        RECT 132.025 69.315 132.195 69.485 ;
        RECT 132.485 69.315 132.655 69.485 ;
        RECT 132.945 69.315 133.115 69.485 ;
        RECT 133.405 69.315 133.575 69.485 ;
        RECT 133.865 69.315 134.035 69.485 ;
        RECT 134.325 69.315 134.495 69.485 ;
        RECT 134.785 69.315 134.955 69.485 ;
        RECT 135.245 69.315 135.415 69.485 ;
        RECT 135.705 69.315 135.875 69.485 ;
        RECT 136.165 69.315 136.335 69.485 ;
        RECT 136.625 69.315 136.795 69.485 ;
        RECT 137.085 69.315 137.255 69.485 ;
        RECT 137.545 69.315 137.715 69.485 ;
        RECT 138.005 69.315 138.175 69.485 ;
        RECT 138.465 69.315 138.635 69.485 ;
        RECT 138.925 69.315 139.095 69.485 ;
        RECT 139.385 69.315 139.555 69.485 ;
        RECT 139.845 69.315 140.015 69.485 ;
        RECT 140.305 69.315 140.475 69.485 ;
        RECT 140.765 69.315 140.935 69.485 ;
        RECT 141.225 69.315 141.395 69.485 ;
        RECT 141.685 69.315 141.855 69.485 ;
        RECT 142.145 69.315 142.315 69.485 ;
        RECT 142.605 69.315 142.775 69.485 ;
        RECT 143.065 69.315 143.235 69.485 ;
        RECT 143.525 69.315 143.695 69.485 ;
        RECT 143.985 69.315 144.155 69.485 ;
        RECT 55.665 63.875 55.835 64.045 ;
        RECT 56.125 63.875 56.295 64.045 ;
        RECT 56.585 63.875 56.755 64.045 ;
        RECT 57.045 63.875 57.215 64.045 ;
        RECT 57.505 63.875 57.675 64.045 ;
        RECT 57.965 63.875 58.135 64.045 ;
        RECT 58.425 63.875 58.595 64.045 ;
        RECT 58.885 63.875 59.055 64.045 ;
        RECT 59.345 63.875 59.515 64.045 ;
        RECT 59.805 63.875 59.975 64.045 ;
        RECT 60.265 63.875 60.435 64.045 ;
        RECT 60.725 63.875 60.895 64.045 ;
        RECT 61.185 63.875 61.355 64.045 ;
        RECT 61.645 63.875 61.815 64.045 ;
        RECT 62.105 63.875 62.275 64.045 ;
        RECT 62.565 63.875 62.735 64.045 ;
        RECT 63.025 63.875 63.195 64.045 ;
        RECT 63.485 63.875 63.655 64.045 ;
        RECT 63.945 63.875 64.115 64.045 ;
        RECT 64.405 63.875 64.575 64.045 ;
        RECT 64.865 63.875 65.035 64.045 ;
        RECT 65.325 63.875 65.495 64.045 ;
        RECT 65.785 63.875 65.955 64.045 ;
        RECT 66.245 63.875 66.415 64.045 ;
        RECT 66.705 63.875 66.875 64.045 ;
        RECT 67.165 63.875 67.335 64.045 ;
        RECT 67.625 63.875 67.795 64.045 ;
        RECT 68.085 63.875 68.255 64.045 ;
        RECT 68.545 63.875 68.715 64.045 ;
        RECT 69.005 63.875 69.175 64.045 ;
        RECT 69.465 63.875 69.635 64.045 ;
        RECT 69.925 63.875 70.095 64.045 ;
        RECT 70.385 63.875 70.555 64.045 ;
        RECT 70.845 63.875 71.015 64.045 ;
        RECT 71.305 63.875 71.475 64.045 ;
        RECT 71.765 63.875 71.935 64.045 ;
        RECT 72.225 63.875 72.395 64.045 ;
        RECT 72.685 63.875 72.855 64.045 ;
        RECT 73.145 63.875 73.315 64.045 ;
        RECT 73.605 63.875 73.775 64.045 ;
        RECT 74.065 63.875 74.235 64.045 ;
        RECT 74.525 63.875 74.695 64.045 ;
        RECT 74.985 63.875 75.155 64.045 ;
        RECT 75.445 63.875 75.615 64.045 ;
        RECT 75.905 63.875 76.075 64.045 ;
        RECT 76.365 63.875 76.535 64.045 ;
        RECT 76.825 63.875 76.995 64.045 ;
        RECT 77.285 63.875 77.455 64.045 ;
        RECT 77.745 63.875 77.915 64.045 ;
        RECT 78.205 63.875 78.375 64.045 ;
        RECT 78.665 63.875 78.835 64.045 ;
        RECT 79.125 63.875 79.295 64.045 ;
        RECT 79.585 63.875 79.755 64.045 ;
        RECT 80.045 63.875 80.215 64.045 ;
        RECT 80.505 63.875 80.675 64.045 ;
        RECT 80.965 63.875 81.135 64.045 ;
        RECT 81.425 63.875 81.595 64.045 ;
        RECT 81.885 63.875 82.055 64.045 ;
        RECT 82.345 63.875 82.515 64.045 ;
        RECT 82.805 63.875 82.975 64.045 ;
        RECT 83.265 63.875 83.435 64.045 ;
        RECT 83.725 63.875 83.895 64.045 ;
        RECT 84.185 63.875 84.355 64.045 ;
        RECT 84.645 63.875 84.815 64.045 ;
        RECT 85.105 63.875 85.275 64.045 ;
        RECT 85.565 63.875 85.735 64.045 ;
        RECT 86.025 63.875 86.195 64.045 ;
        RECT 86.485 63.875 86.655 64.045 ;
        RECT 86.945 63.875 87.115 64.045 ;
        RECT 87.405 63.875 87.575 64.045 ;
        RECT 87.865 63.875 88.035 64.045 ;
        RECT 88.325 63.875 88.495 64.045 ;
        RECT 88.785 63.875 88.955 64.045 ;
        RECT 89.245 63.875 89.415 64.045 ;
        RECT 89.705 63.875 89.875 64.045 ;
        RECT 90.165 63.875 90.335 64.045 ;
        RECT 90.625 63.875 90.795 64.045 ;
        RECT 91.085 63.875 91.255 64.045 ;
        RECT 91.545 63.875 91.715 64.045 ;
        RECT 92.005 63.875 92.175 64.045 ;
        RECT 92.465 63.875 92.635 64.045 ;
        RECT 92.925 63.875 93.095 64.045 ;
        RECT 93.385 63.875 93.555 64.045 ;
        RECT 93.845 63.875 94.015 64.045 ;
        RECT 94.305 63.875 94.475 64.045 ;
        RECT 94.765 63.875 94.935 64.045 ;
        RECT 95.225 63.875 95.395 64.045 ;
        RECT 95.685 63.875 95.855 64.045 ;
        RECT 96.145 63.875 96.315 64.045 ;
        RECT 96.605 63.875 96.775 64.045 ;
        RECT 97.065 63.875 97.235 64.045 ;
        RECT 97.525 63.875 97.695 64.045 ;
        RECT 97.985 63.875 98.155 64.045 ;
        RECT 98.445 63.875 98.615 64.045 ;
        RECT 98.905 63.875 99.075 64.045 ;
        RECT 99.365 63.875 99.535 64.045 ;
        RECT 99.825 63.875 99.995 64.045 ;
        RECT 100.285 63.875 100.455 64.045 ;
        RECT 100.745 63.875 100.915 64.045 ;
        RECT 101.205 63.875 101.375 64.045 ;
        RECT 101.665 63.875 101.835 64.045 ;
        RECT 102.125 63.875 102.295 64.045 ;
        RECT 102.585 63.875 102.755 64.045 ;
        RECT 103.045 63.875 103.215 64.045 ;
        RECT 103.505 63.875 103.675 64.045 ;
        RECT 103.965 63.875 104.135 64.045 ;
        RECT 104.425 63.875 104.595 64.045 ;
        RECT 104.885 63.875 105.055 64.045 ;
        RECT 105.345 63.875 105.515 64.045 ;
        RECT 105.805 63.875 105.975 64.045 ;
        RECT 106.265 63.875 106.435 64.045 ;
        RECT 106.725 63.875 106.895 64.045 ;
        RECT 107.185 63.875 107.355 64.045 ;
        RECT 107.645 63.875 107.815 64.045 ;
        RECT 108.105 63.875 108.275 64.045 ;
        RECT 108.565 63.875 108.735 64.045 ;
        RECT 109.025 63.875 109.195 64.045 ;
        RECT 109.485 63.875 109.655 64.045 ;
        RECT 109.945 63.875 110.115 64.045 ;
        RECT 110.405 63.875 110.575 64.045 ;
        RECT 110.865 63.875 111.035 64.045 ;
        RECT 111.325 63.875 111.495 64.045 ;
        RECT 111.785 63.875 111.955 64.045 ;
        RECT 112.245 63.875 112.415 64.045 ;
        RECT 112.705 63.875 112.875 64.045 ;
        RECT 113.165 63.875 113.335 64.045 ;
        RECT 113.625 63.875 113.795 64.045 ;
        RECT 114.085 63.875 114.255 64.045 ;
        RECT 114.545 63.875 114.715 64.045 ;
        RECT 115.005 63.875 115.175 64.045 ;
        RECT 115.465 63.875 115.635 64.045 ;
        RECT 115.925 63.875 116.095 64.045 ;
        RECT 116.385 63.875 116.555 64.045 ;
        RECT 116.845 63.875 117.015 64.045 ;
        RECT 117.305 63.875 117.475 64.045 ;
        RECT 117.765 63.875 117.935 64.045 ;
        RECT 118.225 63.875 118.395 64.045 ;
        RECT 118.685 63.875 118.855 64.045 ;
        RECT 119.145 63.875 119.315 64.045 ;
        RECT 119.605 63.875 119.775 64.045 ;
        RECT 120.065 63.875 120.235 64.045 ;
        RECT 120.525 63.875 120.695 64.045 ;
        RECT 120.985 63.875 121.155 64.045 ;
        RECT 121.445 63.875 121.615 64.045 ;
        RECT 121.905 63.875 122.075 64.045 ;
        RECT 122.365 63.875 122.535 64.045 ;
        RECT 122.825 63.875 122.995 64.045 ;
        RECT 123.285 63.875 123.455 64.045 ;
        RECT 123.745 63.875 123.915 64.045 ;
        RECT 124.205 63.875 124.375 64.045 ;
        RECT 124.665 63.875 124.835 64.045 ;
        RECT 125.125 63.875 125.295 64.045 ;
        RECT 125.585 63.875 125.755 64.045 ;
        RECT 126.045 63.875 126.215 64.045 ;
        RECT 126.505 63.875 126.675 64.045 ;
        RECT 126.965 63.875 127.135 64.045 ;
        RECT 127.425 63.875 127.595 64.045 ;
        RECT 127.885 63.875 128.055 64.045 ;
        RECT 128.345 63.875 128.515 64.045 ;
        RECT 128.805 63.875 128.975 64.045 ;
        RECT 129.265 63.875 129.435 64.045 ;
        RECT 129.725 63.875 129.895 64.045 ;
        RECT 130.185 63.875 130.355 64.045 ;
        RECT 130.645 63.875 130.815 64.045 ;
        RECT 131.105 63.875 131.275 64.045 ;
        RECT 131.565 63.875 131.735 64.045 ;
        RECT 132.025 63.875 132.195 64.045 ;
        RECT 132.485 63.875 132.655 64.045 ;
        RECT 132.945 63.875 133.115 64.045 ;
        RECT 133.405 63.875 133.575 64.045 ;
        RECT 133.865 63.875 134.035 64.045 ;
        RECT 134.325 63.875 134.495 64.045 ;
        RECT 134.785 63.875 134.955 64.045 ;
        RECT 135.245 63.875 135.415 64.045 ;
        RECT 135.705 63.875 135.875 64.045 ;
        RECT 136.165 63.875 136.335 64.045 ;
        RECT 136.625 63.875 136.795 64.045 ;
        RECT 137.085 63.875 137.255 64.045 ;
        RECT 137.545 63.875 137.715 64.045 ;
        RECT 138.005 63.875 138.175 64.045 ;
        RECT 138.465 63.875 138.635 64.045 ;
        RECT 138.925 63.875 139.095 64.045 ;
        RECT 139.385 63.875 139.555 64.045 ;
        RECT 139.845 63.875 140.015 64.045 ;
        RECT 140.305 63.875 140.475 64.045 ;
        RECT 140.765 63.875 140.935 64.045 ;
        RECT 141.225 63.875 141.395 64.045 ;
        RECT 141.685 63.875 141.855 64.045 ;
        RECT 142.145 63.875 142.315 64.045 ;
        RECT 142.605 63.875 142.775 64.045 ;
        RECT 143.065 63.875 143.235 64.045 ;
        RECT 143.525 63.875 143.695 64.045 ;
        RECT 143.985 63.875 144.155 64.045 ;
        RECT 55.665 58.435 55.835 58.605 ;
        RECT 56.125 58.435 56.295 58.605 ;
        RECT 56.585 58.435 56.755 58.605 ;
        RECT 57.045 58.435 57.215 58.605 ;
        RECT 57.505 58.435 57.675 58.605 ;
        RECT 57.965 58.435 58.135 58.605 ;
        RECT 58.425 58.435 58.595 58.605 ;
        RECT 58.885 58.435 59.055 58.605 ;
        RECT 59.345 58.435 59.515 58.605 ;
        RECT 59.805 58.435 59.975 58.605 ;
        RECT 60.265 58.435 60.435 58.605 ;
        RECT 60.725 58.435 60.895 58.605 ;
        RECT 61.185 58.435 61.355 58.605 ;
        RECT 61.645 58.435 61.815 58.605 ;
        RECT 62.105 58.435 62.275 58.605 ;
        RECT 62.565 58.435 62.735 58.605 ;
        RECT 63.025 58.435 63.195 58.605 ;
        RECT 63.485 58.435 63.655 58.605 ;
        RECT 63.945 58.435 64.115 58.605 ;
        RECT 64.405 58.435 64.575 58.605 ;
        RECT 64.865 58.435 65.035 58.605 ;
        RECT 65.325 58.435 65.495 58.605 ;
        RECT 65.785 58.435 65.955 58.605 ;
        RECT 66.245 58.435 66.415 58.605 ;
        RECT 66.705 58.435 66.875 58.605 ;
        RECT 67.165 58.435 67.335 58.605 ;
        RECT 67.625 58.435 67.795 58.605 ;
        RECT 68.085 58.435 68.255 58.605 ;
        RECT 68.545 58.435 68.715 58.605 ;
        RECT 69.005 58.435 69.175 58.605 ;
        RECT 69.465 58.435 69.635 58.605 ;
        RECT 69.925 58.435 70.095 58.605 ;
        RECT 70.385 58.435 70.555 58.605 ;
        RECT 70.845 58.435 71.015 58.605 ;
        RECT 71.305 58.435 71.475 58.605 ;
        RECT 71.765 58.435 71.935 58.605 ;
        RECT 72.225 58.435 72.395 58.605 ;
        RECT 72.685 58.435 72.855 58.605 ;
        RECT 73.145 58.435 73.315 58.605 ;
        RECT 73.605 58.435 73.775 58.605 ;
        RECT 74.065 58.435 74.235 58.605 ;
        RECT 74.525 58.435 74.695 58.605 ;
        RECT 74.985 58.435 75.155 58.605 ;
        RECT 75.445 58.435 75.615 58.605 ;
        RECT 75.905 58.435 76.075 58.605 ;
        RECT 76.365 58.435 76.535 58.605 ;
        RECT 76.825 58.435 76.995 58.605 ;
        RECT 77.285 58.435 77.455 58.605 ;
        RECT 77.745 58.435 77.915 58.605 ;
        RECT 78.205 58.435 78.375 58.605 ;
        RECT 78.665 58.435 78.835 58.605 ;
        RECT 79.125 58.435 79.295 58.605 ;
        RECT 79.585 58.435 79.755 58.605 ;
        RECT 80.045 58.435 80.215 58.605 ;
        RECT 80.505 58.435 80.675 58.605 ;
        RECT 80.965 58.435 81.135 58.605 ;
        RECT 81.425 58.435 81.595 58.605 ;
        RECT 81.885 58.435 82.055 58.605 ;
        RECT 82.345 58.435 82.515 58.605 ;
        RECT 82.805 58.435 82.975 58.605 ;
        RECT 83.265 58.435 83.435 58.605 ;
        RECT 83.725 58.435 83.895 58.605 ;
        RECT 84.185 58.435 84.355 58.605 ;
        RECT 84.645 58.435 84.815 58.605 ;
        RECT 85.105 58.435 85.275 58.605 ;
        RECT 85.565 58.435 85.735 58.605 ;
        RECT 86.025 58.435 86.195 58.605 ;
        RECT 86.485 58.435 86.655 58.605 ;
        RECT 86.945 58.435 87.115 58.605 ;
        RECT 87.405 58.435 87.575 58.605 ;
        RECT 87.865 58.435 88.035 58.605 ;
        RECT 88.325 58.435 88.495 58.605 ;
        RECT 88.785 58.435 88.955 58.605 ;
        RECT 89.245 58.435 89.415 58.605 ;
        RECT 89.705 58.435 89.875 58.605 ;
        RECT 90.165 58.435 90.335 58.605 ;
        RECT 90.625 58.435 90.795 58.605 ;
        RECT 91.085 58.435 91.255 58.605 ;
        RECT 91.545 58.435 91.715 58.605 ;
        RECT 92.005 58.435 92.175 58.605 ;
        RECT 92.465 58.435 92.635 58.605 ;
        RECT 92.925 58.435 93.095 58.605 ;
        RECT 93.385 58.435 93.555 58.605 ;
        RECT 93.845 58.435 94.015 58.605 ;
        RECT 94.305 58.435 94.475 58.605 ;
        RECT 94.765 58.435 94.935 58.605 ;
        RECT 95.225 58.435 95.395 58.605 ;
        RECT 95.685 58.435 95.855 58.605 ;
        RECT 96.145 58.435 96.315 58.605 ;
        RECT 96.605 58.435 96.775 58.605 ;
        RECT 97.065 58.435 97.235 58.605 ;
        RECT 97.525 58.435 97.695 58.605 ;
        RECT 97.985 58.435 98.155 58.605 ;
        RECT 98.445 58.435 98.615 58.605 ;
        RECT 98.905 58.435 99.075 58.605 ;
        RECT 99.365 58.435 99.535 58.605 ;
        RECT 99.825 58.435 99.995 58.605 ;
        RECT 100.285 58.435 100.455 58.605 ;
        RECT 100.745 58.435 100.915 58.605 ;
        RECT 101.205 58.435 101.375 58.605 ;
        RECT 101.665 58.435 101.835 58.605 ;
        RECT 102.125 58.435 102.295 58.605 ;
        RECT 102.585 58.435 102.755 58.605 ;
        RECT 103.045 58.435 103.215 58.605 ;
        RECT 103.505 58.435 103.675 58.605 ;
        RECT 103.965 58.435 104.135 58.605 ;
        RECT 104.425 58.435 104.595 58.605 ;
        RECT 104.885 58.435 105.055 58.605 ;
        RECT 105.345 58.435 105.515 58.605 ;
        RECT 105.805 58.435 105.975 58.605 ;
        RECT 106.265 58.435 106.435 58.605 ;
        RECT 106.725 58.435 106.895 58.605 ;
        RECT 107.185 58.435 107.355 58.605 ;
        RECT 107.645 58.435 107.815 58.605 ;
        RECT 108.105 58.435 108.275 58.605 ;
        RECT 108.565 58.435 108.735 58.605 ;
        RECT 109.025 58.435 109.195 58.605 ;
        RECT 109.485 58.435 109.655 58.605 ;
        RECT 109.945 58.435 110.115 58.605 ;
        RECT 110.405 58.435 110.575 58.605 ;
        RECT 110.865 58.435 111.035 58.605 ;
        RECT 111.325 58.435 111.495 58.605 ;
        RECT 111.785 58.435 111.955 58.605 ;
        RECT 112.245 58.435 112.415 58.605 ;
        RECT 112.705 58.435 112.875 58.605 ;
        RECT 113.165 58.435 113.335 58.605 ;
        RECT 113.625 58.435 113.795 58.605 ;
        RECT 114.085 58.435 114.255 58.605 ;
        RECT 114.545 58.435 114.715 58.605 ;
        RECT 115.005 58.435 115.175 58.605 ;
        RECT 115.465 58.435 115.635 58.605 ;
        RECT 115.925 58.435 116.095 58.605 ;
        RECT 116.385 58.435 116.555 58.605 ;
        RECT 116.845 58.435 117.015 58.605 ;
        RECT 117.305 58.435 117.475 58.605 ;
        RECT 117.765 58.435 117.935 58.605 ;
        RECT 118.225 58.435 118.395 58.605 ;
        RECT 118.685 58.435 118.855 58.605 ;
        RECT 119.145 58.435 119.315 58.605 ;
        RECT 119.605 58.435 119.775 58.605 ;
        RECT 120.065 58.435 120.235 58.605 ;
        RECT 120.525 58.435 120.695 58.605 ;
        RECT 120.985 58.435 121.155 58.605 ;
        RECT 121.445 58.435 121.615 58.605 ;
        RECT 121.905 58.435 122.075 58.605 ;
        RECT 122.365 58.435 122.535 58.605 ;
        RECT 122.825 58.435 122.995 58.605 ;
        RECT 123.285 58.435 123.455 58.605 ;
        RECT 123.745 58.435 123.915 58.605 ;
        RECT 124.205 58.435 124.375 58.605 ;
        RECT 124.665 58.435 124.835 58.605 ;
        RECT 125.125 58.435 125.295 58.605 ;
        RECT 125.585 58.435 125.755 58.605 ;
        RECT 126.045 58.435 126.215 58.605 ;
        RECT 126.505 58.435 126.675 58.605 ;
        RECT 126.965 58.435 127.135 58.605 ;
        RECT 127.425 58.435 127.595 58.605 ;
        RECT 127.885 58.435 128.055 58.605 ;
        RECT 128.345 58.435 128.515 58.605 ;
        RECT 128.805 58.435 128.975 58.605 ;
        RECT 129.265 58.435 129.435 58.605 ;
        RECT 129.725 58.435 129.895 58.605 ;
        RECT 130.185 58.435 130.355 58.605 ;
        RECT 130.645 58.435 130.815 58.605 ;
        RECT 131.105 58.435 131.275 58.605 ;
        RECT 131.565 58.435 131.735 58.605 ;
        RECT 132.025 58.435 132.195 58.605 ;
        RECT 132.485 58.435 132.655 58.605 ;
        RECT 132.945 58.435 133.115 58.605 ;
        RECT 133.405 58.435 133.575 58.605 ;
        RECT 133.865 58.435 134.035 58.605 ;
        RECT 134.325 58.435 134.495 58.605 ;
        RECT 134.785 58.435 134.955 58.605 ;
        RECT 135.245 58.435 135.415 58.605 ;
        RECT 135.705 58.435 135.875 58.605 ;
        RECT 136.165 58.435 136.335 58.605 ;
        RECT 136.625 58.435 136.795 58.605 ;
        RECT 137.085 58.435 137.255 58.605 ;
        RECT 137.545 58.435 137.715 58.605 ;
        RECT 138.005 58.435 138.175 58.605 ;
        RECT 138.465 58.435 138.635 58.605 ;
        RECT 138.925 58.435 139.095 58.605 ;
        RECT 139.385 58.435 139.555 58.605 ;
        RECT 139.845 58.435 140.015 58.605 ;
        RECT 140.305 58.435 140.475 58.605 ;
        RECT 140.765 58.435 140.935 58.605 ;
        RECT 141.225 58.435 141.395 58.605 ;
        RECT 141.685 58.435 141.855 58.605 ;
        RECT 142.145 58.435 142.315 58.605 ;
        RECT 142.605 58.435 142.775 58.605 ;
        RECT 143.065 58.435 143.235 58.605 ;
        RECT 143.525 58.435 143.695 58.605 ;
        RECT 143.985 58.435 144.155 58.605 ;
        RECT 55.665 52.995 55.835 53.165 ;
        RECT 56.125 52.995 56.295 53.165 ;
        RECT 56.585 52.995 56.755 53.165 ;
        RECT 57.045 52.995 57.215 53.165 ;
        RECT 57.505 52.995 57.675 53.165 ;
        RECT 57.965 52.995 58.135 53.165 ;
        RECT 58.425 52.995 58.595 53.165 ;
        RECT 58.885 52.995 59.055 53.165 ;
        RECT 59.345 52.995 59.515 53.165 ;
        RECT 59.805 52.995 59.975 53.165 ;
        RECT 60.265 52.995 60.435 53.165 ;
        RECT 60.725 52.995 60.895 53.165 ;
        RECT 61.185 52.995 61.355 53.165 ;
        RECT 61.645 52.995 61.815 53.165 ;
        RECT 62.105 52.995 62.275 53.165 ;
        RECT 62.565 52.995 62.735 53.165 ;
        RECT 63.025 52.995 63.195 53.165 ;
        RECT 63.485 52.995 63.655 53.165 ;
        RECT 63.945 52.995 64.115 53.165 ;
        RECT 64.405 52.995 64.575 53.165 ;
        RECT 64.865 52.995 65.035 53.165 ;
        RECT 65.325 52.995 65.495 53.165 ;
        RECT 65.785 52.995 65.955 53.165 ;
        RECT 66.245 52.995 66.415 53.165 ;
        RECT 66.705 52.995 66.875 53.165 ;
        RECT 67.165 52.995 67.335 53.165 ;
        RECT 67.625 52.995 67.795 53.165 ;
        RECT 68.085 52.995 68.255 53.165 ;
        RECT 68.545 52.995 68.715 53.165 ;
        RECT 69.005 52.995 69.175 53.165 ;
        RECT 69.465 52.995 69.635 53.165 ;
        RECT 69.925 52.995 70.095 53.165 ;
        RECT 70.385 52.995 70.555 53.165 ;
        RECT 70.845 52.995 71.015 53.165 ;
        RECT 71.305 52.995 71.475 53.165 ;
        RECT 71.765 52.995 71.935 53.165 ;
        RECT 72.225 52.995 72.395 53.165 ;
        RECT 72.685 52.995 72.855 53.165 ;
        RECT 73.145 52.995 73.315 53.165 ;
        RECT 73.605 52.995 73.775 53.165 ;
        RECT 74.065 52.995 74.235 53.165 ;
        RECT 74.525 52.995 74.695 53.165 ;
        RECT 74.985 52.995 75.155 53.165 ;
        RECT 75.445 52.995 75.615 53.165 ;
        RECT 75.905 52.995 76.075 53.165 ;
        RECT 76.365 52.995 76.535 53.165 ;
        RECT 76.825 52.995 76.995 53.165 ;
        RECT 77.285 52.995 77.455 53.165 ;
        RECT 77.745 52.995 77.915 53.165 ;
        RECT 78.205 52.995 78.375 53.165 ;
        RECT 78.665 52.995 78.835 53.165 ;
        RECT 79.125 52.995 79.295 53.165 ;
        RECT 79.585 52.995 79.755 53.165 ;
        RECT 80.045 52.995 80.215 53.165 ;
        RECT 80.505 52.995 80.675 53.165 ;
        RECT 80.965 52.995 81.135 53.165 ;
        RECT 81.425 52.995 81.595 53.165 ;
        RECT 81.885 52.995 82.055 53.165 ;
        RECT 82.345 52.995 82.515 53.165 ;
        RECT 82.805 52.995 82.975 53.165 ;
        RECT 83.265 52.995 83.435 53.165 ;
        RECT 83.725 52.995 83.895 53.165 ;
        RECT 84.185 52.995 84.355 53.165 ;
        RECT 84.645 52.995 84.815 53.165 ;
        RECT 85.105 52.995 85.275 53.165 ;
        RECT 85.565 52.995 85.735 53.165 ;
        RECT 86.025 52.995 86.195 53.165 ;
        RECT 86.485 52.995 86.655 53.165 ;
        RECT 86.945 52.995 87.115 53.165 ;
        RECT 87.405 52.995 87.575 53.165 ;
        RECT 87.865 52.995 88.035 53.165 ;
        RECT 88.325 52.995 88.495 53.165 ;
        RECT 88.785 52.995 88.955 53.165 ;
        RECT 89.245 52.995 89.415 53.165 ;
        RECT 89.705 52.995 89.875 53.165 ;
        RECT 90.165 52.995 90.335 53.165 ;
        RECT 90.625 52.995 90.795 53.165 ;
        RECT 91.085 52.995 91.255 53.165 ;
        RECT 91.545 52.995 91.715 53.165 ;
        RECT 92.005 52.995 92.175 53.165 ;
        RECT 92.465 52.995 92.635 53.165 ;
        RECT 92.925 52.995 93.095 53.165 ;
        RECT 93.385 52.995 93.555 53.165 ;
        RECT 93.845 52.995 94.015 53.165 ;
        RECT 94.305 52.995 94.475 53.165 ;
        RECT 94.765 52.995 94.935 53.165 ;
        RECT 95.225 52.995 95.395 53.165 ;
        RECT 95.685 52.995 95.855 53.165 ;
        RECT 96.145 52.995 96.315 53.165 ;
        RECT 96.605 52.995 96.775 53.165 ;
        RECT 97.065 52.995 97.235 53.165 ;
        RECT 97.525 52.995 97.695 53.165 ;
        RECT 97.985 52.995 98.155 53.165 ;
        RECT 98.445 52.995 98.615 53.165 ;
        RECT 98.905 52.995 99.075 53.165 ;
        RECT 99.365 52.995 99.535 53.165 ;
        RECT 99.825 52.995 99.995 53.165 ;
        RECT 100.285 52.995 100.455 53.165 ;
        RECT 100.745 52.995 100.915 53.165 ;
        RECT 101.205 52.995 101.375 53.165 ;
        RECT 101.665 52.995 101.835 53.165 ;
        RECT 102.125 52.995 102.295 53.165 ;
        RECT 102.585 52.995 102.755 53.165 ;
        RECT 103.045 52.995 103.215 53.165 ;
        RECT 103.505 52.995 103.675 53.165 ;
        RECT 103.965 52.995 104.135 53.165 ;
        RECT 104.425 52.995 104.595 53.165 ;
        RECT 104.885 52.995 105.055 53.165 ;
        RECT 105.345 52.995 105.515 53.165 ;
        RECT 105.805 52.995 105.975 53.165 ;
        RECT 106.265 52.995 106.435 53.165 ;
        RECT 106.725 52.995 106.895 53.165 ;
        RECT 107.185 52.995 107.355 53.165 ;
        RECT 107.645 52.995 107.815 53.165 ;
        RECT 108.105 52.995 108.275 53.165 ;
        RECT 108.565 52.995 108.735 53.165 ;
        RECT 109.025 52.995 109.195 53.165 ;
        RECT 109.485 52.995 109.655 53.165 ;
        RECT 109.945 52.995 110.115 53.165 ;
        RECT 110.405 52.995 110.575 53.165 ;
        RECT 110.865 52.995 111.035 53.165 ;
        RECT 111.325 52.995 111.495 53.165 ;
        RECT 111.785 52.995 111.955 53.165 ;
        RECT 112.245 52.995 112.415 53.165 ;
        RECT 112.705 52.995 112.875 53.165 ;
        RECT 113.165 52.995 113.335 53.165 ;
        RECT 113.625 52.995 113.795 53.165 ;
        RECT 114.085 52.995 114.255 53.165 ;
        RECT 114.545 52.995 114.715 53.165 ;
        RECT 115.005 52.995 115.175 53.165 ;
        RECT 115.465 52.995 115.635 53.165 ;
        RECT 115.925 52.995 116.095 53.165 ;
        RECT 116.385 52.995 116.555 53.165 ;
        RECT 116.845 52.995 117.015 53.165 ;
        RECT 117.305 52.995 117.475 53.165 ;
        RECT 117.765 52.995 117.935 53.165 ;
        RECT 118.225 52.995 118.395 53.165 ;
        RECT 118.685 52.995 118.855 53.165 ;
        RECT 119.145 52.995 119.315 53.165 ;
        RECT 119.605 52.995 119.775 53.165 ;
        RECT 120.065 52.995 120.235 53.165 ;
        RECT 120.525 52.995 120.695 53.165 ;
        RECT 120.985 52.995 121.155 53.165 ;
        RECT 121.445 52.995 121.615 53.165 ;
        RECT 121.905 52.995 122.075 53.165 ;
        RECT 122.365 52.995 122.535 53.165 ;
        RECT 122.825 52.995 122.995 53.165 ;
        RECT 123.285 52.995 123.455 53.165 ;
        RECT 123.745 52.995 123.915 53.165 ;
        RECT 124.205 52.995 124.375 53.165 ;
        RECT 124.665 52.995 124.835 53.165 ;
        RECT 125.125 52.995 125.295 53.165 ;
        RECT 125.585 52.995 125.755 53.165 ;
        RECT 126.045 52.995 126.215 53.165 ;
        RECT 126.505 52.995 126.675 53.165 ;
        RECT 126.965 52.995 127.135 53.165 ;
        RECT 127.425 52.995 127.595 53.165 ;
        RECT 127.885 52.995 128.055 53.165 ;
        RECT 128.345 52.995 128.515 53.165 ;
        RECT 128.805 52.995 128.975 53.165 ;
        RECT 129.265 52.995 129.435 53.165 ;
        RECT 129.725 52.995 129.895 53.165 ;
        RECT 130.185 52.995 130.355 53.165 ;
        RECT 130.645 52.995 130.815 53.165 ;
        RECT 131.105 52.995 131.275 53.165 ;
        RECT 131.565 52.995 131.735 53.165 ;
        RECT 132.025 52.995 132.195 53.165 ;
        RECT 132.485 52.995 132.655 53.165 ;
        RECT 132.945 52.995 133.115 53.165 ;
        RECT 133.405 52.995 133.575 53.165 ;
        RECT 133.865 52.995 134.035 53.165 ;
        RECT 134.325 52.995 134.495 53.165 ;
        RECT 134.785 52.995 134.955 53.165 ;
        RECT 135.245 52.995 135.415 53.165 ;
        RECT 135.705 52.995 135.875 53.165 ;
        RECT 136.165 52.995 136.335 53.165 ;
        RECT 136.625 52.995 136.795 53.165 ;
        RECT 137.085 52.995 137.255 53.165 ;
        RECT 137.545 52.995 137.715 53.165 ;
        RECT 138.005 52.995 138.175 53.165 ;
        RECT 138.465 52.995 138.635 53.165 ;
        RECT 138.925 52.995 139.095 53.165 ;
        RECT 139.385 52.995 139.555 53.165 ;
        RECT 139.845 52.995 140.015 53.165 ;
        RECT 140.305 52.995 140.475 53.165 ;
        RECT 140.765 52.995 140.935 53.165 ;
        RECT 141.225 52.995 141.395 53.165 ;
        RECT 141.685 52.995 141.855 53.165 ;
        RECT 142.145 52.995 142.315 53.165 ;
        RECT 142.605 52.995 142.775 53.165 ;
        RECT 143.065 52.995 143.235 53.165 ;
        RECT 143.525 52.995 143.695 53.165 ;
        RECT 143.985 52.995 144.155 53.165 ;
        RECT 55.665 47.555 55.835 47.725 ;
        RECT 56.125 47.555 56.295 47.725 ;
        RECT 56.585 47.555 56.755 47.725 ;
        RECT 57.045 47.555 57.215 47.725 ;
        RECT 57.505 47.555 57.675 47.725 ;
        RECT 57.965 47.555 58.135 47.725 ;
        RECT 58.425 47.555 58.595 47.725 ;
        RECT 58.885 47.555 59.055 47.725 ;
        RECT 59.345 47.555 59.515 47.725 ;
        RECT 59.805 47.555 59.975 47.725 ;
        RECT 60.265 47.555 60.435 47.725 ;
        RECT 60.725 47.555 60.895 47.725 ;
        RECT 61.185 47.555 61.355 47.725 ;
        RECT 61.645 47.555 61.815 47.725 ;
        RECT 62.105 47.555 62.275 47.725 ;
        RECT 62.565 47.555 62.735 47.725 ;
        RECT 63.025 47.555 63.195 47.725 ;
        RECT 63.485 47.555 63.655 47.725 ;
        RECT 63.945 47.555 64.115 47.725 ;
        RECT 64.405 47.555 64.575 47.725 ;
        RECT 64.865 47.555 65.035 47.725 ;
        RECT 65.325 47.555 65.495 47.725 ;
        RECT 65.785 47.555 65.955 47.725 ;
        RECT 66.245 47.555 66.415 47.725 ;
        RECT 66.705 47.555 66.875 47.725 ;
        RECT 67.165 47.555 67.335 47.725 ;
        RECT 67.625 47.555 67.795 47.725 ;
        RECT 68.085 47.555 68.255 47.725 ;
        RECT 68.545 47.555 68.715 47.725 ;
        RECT 69.005 47.555 69.175 47.725 ;
        RECT 69.465 47.555 69.635 47.725 ;
        RECT 69.925 47.555 70.095 47.725 ;
        RECT 70.385 47.555 70.555 47.725 ;
        RECT 70.845 47.555 71.015 47.725 ;
        RECT 71.305 47.555 71.475 47.725 ;
        RECT 71.765 47.555 71.935 47.725 ;
        RECT 72.225 47.555 72.395 47.725 ;
        RECT 72.685 47.555 72.855 47.725 ;
        RECT 73.145 47.555 73.315 47.725 ;
        RECT 73.605 47.555 73.775 47.725 ;
        RECT 74.065 47.555 74.235 47.725 ;
        RECT 74.525 47.555 74.695 47.725 ;
        RECT 74.985 47.555 75.155 47.725 ;
        RECT 75.445 47.555 75.615 47.725 ;
        RECT 75.905 47.555 76.075 47.725 ;
        RECT 76.365 47.555 76.535 47.725 ;
        RECT 76.825 47.555 76.995 47.725 ;
        RECT 77.285 47.555 77.455 47.725 ;
        RECT 77.745 47.555 77.915 47.725 ;
        RECT 78.205 47.555 78.375 47.725 ;
        RECT 78.665 47.555 78.835 47.725 ;
        RECT 79.125 47.555 79.295 47.725 ;
        RECT 79.585 47.555 79.755 47.725 ;
        RECT 80.045 47.555 80.215 47.725 ;
        RECT 80.505 47.555 80.675 47.725 ;
        RECT 80.965 47.555 81.135 47.725 ;
        RECT 81.425 47.555 81.595 47.725 ;
        RECT 81.885 47.555 82.055 47.725 ;
        RECT 82.345 47.555 82.515 47.725 ;
        RECT 82.805 47.555 82.975 47.725 ;
        RECT 83.265 47.555 83.435 47.725 ;
        RECT 83.725 47.555 83.895 47.725 ;
        RECT 84.185 47.555 84.355 47.725 ;
        RECT 84.645 47.555 84.815 47.725 ;
        RECT 85.105 47.555 85.275 47.725 ;
        RECT 85.565 47.555 85.735 47.725 ;
        RECT 86.025 47.555 86.195 47.725 ;
        RECT 86.485 47.555 86.655 47.725 ;
        RECT 86.945 47.555 87.115 47.725 ;
        RECT 87.405 47.555 87.575 47.725 ;
        RECT 87.865 47.555 88.035 47.725 ;
        RECT 88.325 47.555 88.495 47.725 ;
        RECT 88.785 47.555 88.955 47.725 ;
        RECT 89.245 47.555 89.415 47.725 ;
        RECT 89.705 47.555 89.875 47.725 ;
        RECT 90.165 47.555 90.335 47.725 ;
        RECT 90.625 47.555 90.795 47.725 ;
        RECT 91.085 47.555 91.255 47.725 ;
        RECT 91.545 47.555 91.715 47.725 ;
        RECT 92.005 47.555 92.175 47.725 ;
        RECT 92.465 47.555 92.635 47.725 ;
        RECT 92.925 47.555 93.095 47.725 ;
        RECT 93.385 47.555 93.555 47.725 ;
        RECT 93.845 47.555 94.015 47.725 ;
        RECT 94.305 47.555 94.475 47.725 ;
        RECT 94.765 47.555 94.935 47.725 ;
        RECT 95.225 47.555 95.395 47.725 ;
        RECT 95.685 47.555 95.855 47.725 ;
        RECT 96.145 47.555 96.315 47.725 ;
        RECT 96.605 47.555 96.775 47.725 ;
        RECT 97.065 47.555 97.235 47.725 ;
        RECT 97.525 47.555 97.695 47.725 ;
        RECT 97.985 47.555 98.155 47.725 ;
        RECT 98.445 47.555 98.615 47.725 ;
        RECT 98.905 47.555 99.075 47.725 ;
        RECT 99.365 47.555 99.535 47.725 ;
        RECT 99.825 47.555 99.995 47.725 ;
        RECT 100.285 47.555 100.455 47.725 ;
        RECT 100.745 47.555 100.915 47.725 ;
        RECT 101.205 47.555 101.375 47.725 ;
        RECT 101.665 47.555 101.835 47.725 ;
        RECT 102.125 47.555 102.295 47.725 ;
        RECT 102.585 47.555 102.755 47.725 ;
        RECT 103.045 47.555 103.215 47.725 ;
        RECT 103.505 47.555 103.675 47.725 ;
        RECT 103.965 47.555 104.135 47.725 ;
        RECT 104.425 47.555 104.595 47.725 ;
        RECT 104.885 47.555 105.055 47.725 ;
        RECT 105.345 47.555 105.515 47.725 ;
        RECT 105.805 47.555 105.975 47.725 ;
        RECT 106.265 47.555 106.435 47.725 ;
        RECT 106.725 47.555 106.895 47.725 ;
        RECT 107.185 47.555 107.355 47.725 ;
        RECT 107.645 47.555 107.815 47.725 ;
        RECT 108.105 47.555 108.275 47.725 ;
        RECT 108.565 47.555 108.735 47.725 ;
        RECT 109.025 47.555 109.195 47.725 ;
        RECT 109.485 47.555 109.655 47.725 ;
        RECT 109.945 47.555 110.115 47.725 ;
        RECT 110.405 47.555 110.575 47.725 ;
        RECT 110.865 47.555 111.035 47.725 ;
        RECT 111.325 47.555 111.495 47.725 ;
        RECT 111.785 47.555 111.955 47.725 ;
        RECT 112.245 47.555 112.415 47.725 ;
        RECT 112.705 47.555 112.875 47.725 ;
        RECT 113.165 47.555 113.335 47.725 ;
        RECT 113.625 47.555 113.795 47.725 ;
        RECT 114.085 47.555 114.255 47.725 ;
        RECT 114.545 47.555 114.715 47.725 ;
        RECT 115.005 47.555 115.175 47.725 ;
        RECT 115.465 47.555 115.635 47.725 ;
        RECT 115.925 47.555 116.095 47.725 ;
        RECT 116.385 47.555 116.555 47.725 ;
        RECT 116.845 47.555 117.015 47.725 ;
        RECT 117.305 47.555 117.475 47.725 ;
        RECT 117.765 47.555 117.935 47.725 ;
        RECT 118.225 47.555 118.395 47.725 ;
        RECT 118.685 47.555 118.855 47.725 ;
        RECT 119.145 47.555 119.315 47.725 ;
        RECT 119.605 47.555 119.775 47.725 ;
        RECT 120.065 47.555 120.235 47.725 ;
        RECT 120.525 47.555 120.695 47.725 ;
        RECT 120.985 47.555 121.155 47.725 ;
        RECT 121.445 47.555 121.615 47.725 ;
        RECT 121.905 47.555 122.075 47.725 ;
        RECT 122.365 47.555 122.535 47.725 ;
        RECT 122.825 47.555 122.995 47.725 ;
        RECT 123.285 47.555 123.455 47.725 ;
        RECT 123.745 47.555 123.915 47.725 ;
        RECT 124.205 47.555 124.375 47.725 ;
        RECT 124.665 47.555 124.835 47.725 ;
        RECT 125.125 47.555 125.295 47.725 ;
        RECT 125.585 47.555 125.755 47.725 ;
        RECT 126.045 47.555 126.215 47.725 ;
        RECT 126.505 47.555 126.675 47.725 ;
        RECT 126.965 47.555 127.135 47.725 ;
        RECT 127.425 47.555 127.595 47.725 ;
        RECT 127.885 47.555 128.055 47.725 ;
        RECT 128.345 47.555 128.515 47.725 ;
        RECT 128.805 47.555 128.975 47.725 ;
        RECT 129.265 47.555 129.435 47.725 ;
        RECT 129.725 47.555 129.895 47.725 ;
        RECT 130.185 47.555 130.355 47.725 ;
        RECT 130.645 47.555 130.815 47.725 ;
        RECT 131.105 47.555 131.275 47.725 ;
        RECT 131.565 47.555 131.735 47.725 ;
        RECT 132.025 47.555 132.195 47.725 ;
        RECT 132.485 47.555 132.655 47.725 ;
        RECT 132.945 47.555 133.115 47.725 ;
        RECT 133.405 47.555 133.575 47.725 ;
        RECT 133.865 47.555 134.035 47.725 ;
        RECT 134.325 47.555 134.495 47.725 ;
        RECT 134.785 47.555 134.955 47.725 ;
        RECT 135.245 47.555 135.415 47.725 ;
        RECT 135.705 47.555 135.875 47.725 ;
        RECT 136.165 47.555 136.335 47.725 ;
        RECT 136.625 47.555 136.795 47.725 ;
        RECT 137.085 47.555 137.255 47.725 ;
        RECT 137.545 47.555 137.715 47.725 ;
        RECT 138.005 47.555 138.175 47.725 ;
        RECT 138.465 47.555 138.635 47.725 ;
        RECT 138.925 47.555 139.095 47.725 ;
        RECT 139.385 47.555 139.555 47.725 ;
        RECT 139.845 47.555 140.015 47.725 ;
        RECT 140.305 47.555 140.475 47.725 ;
        RECT 140.765 47.555 140.935 47.725 ;
        RECT 141.225 47.555 141.395 47.725 ;
        RECT 141.685 47.555 141.855 47.725 ;
        RECT 142.145 47.555 142.315 47.725 ;
        RECT 142.605 47.555 142.775 47.725 ;
        RECT 143.065 47.555 143.235 47.725 ;
        RECT 143.525 47.555 143.695 47.725 ;
        RECT 143.985 47.555 144.155 47.725 ;
        RECT 55.665 42.115 55.835 42.285 ;
        RECT 56.125 42.115 56.295 42.285 ;
        RECT 56.585 42.115 56.755 42.285 ;
        RECT 57.045 42.115 57.215 42.285 ;
        RECT 57.505 42.115 57.675 42.285 ;
        RECT 57.965 42.115 58.135 42.285 ;
        RECT 58.425 42.115 58.595 42.285 ;
        RECT 58.885 42.115 59.055 42.285 ;
        RECT 59.345 42.115 59.515 42.285 ;
        RECT 59.805 42.115 59.975 42.285 ;
        RECT 60.265 42.115 60.435 42.285 ;
        RECT 60.725 42.115 60.895 42.285 ;
        RECT 61.185 42.115 61.355 42.285 ;
        RECT 61.645 42.115 61.815 42.285 ;
        RECT 62.105 42.115 62.275 42.285 ;
        RECT 62.565 42.115 62.735 42.285 ;
        RECT 63.025 42.115 63.195 42.285 ;
        RECT 63.485 42.115 63.655 42.285 ;
        RECT 63.945 42.115 64.115 42.285 ;
        RECT 64.405 42.115 64.575 42.285 ;
        RECT 64.865 42.115 65.035 42.285 ;
        RECT 65.325 42.115 65.495 42.285 ;
        RECT 65.785 42.115 65.955 42.285 ;
        RECT 66.245 42.115 66.415 42.285 ;
        RECT 66.705 42.115 66.875 42.285 ;
        RECT 67.165 42.115 67.335 42.285 ;
        RECT 67.625 42.115 67.795 42.285 ;
        RECT 68.085 42.115 68.255 42.285 ;
        RECT 68.545 42.115 68.715 42.285 ;
        RECT 69.005 42.115 69.175 42.285 ;
        RECT 69.465 42.115 69.635 42.285 ;
        RECT 69.925 42.115 70.095 42.285 ;
        RECT 70.385 42.115 70.555 42.285 ;
        RECT 70.845 42.115 71.015 42.285 ;
        RECT 71.305 42.115 71.475 42.285 ;
        RECT 71.765 42.115 71.935 42.285 ;
        RECT 72.225 42.115 72.395 42.285 ;
        RECT 72.685 42.115 72.855 42.285 ;
        RECT 73.145 42.115 73.315 42.285 ;
        RECT 73.605 42.115 73.775 42.285 ;
        RECT 74.065 42.115 74.235 42.285 ;
        RECT 74.525 42.115 74.695 42.285 ;
        RECT 74.985 42.115 75.155 42.285 ;
        RECT 75.445 42.115 75.615 42.285 ;
        RECT 75.905 42.115 76.075 42.285 ;
        RECT 76.365 42.115 76.535 42.285 ;
        RECT 76.825 42.115 76.995 42.285 ;
        RECT 77.285 42.115 77.455 42.285 ;
        RECT 77.745 42.115 77.915 42.285 ;
        RECT 78.205 42.115 78.375 42.285 ;
        RECT 78.665 42.115 78.835 42.285 ;
        RECT 79.125 42.115 79.295 42.285 ;
        RECT 79.585 42.115 79.755 42.285 ;
        RECT 80.045 42.115 80.215 42.285 ;
        RECT 80.505 42.115 80.675 42.285 ;
        RECT 80.965 42.115 81.135 42.285 ;
        RECT 81.425 42.115 81.595 42.285 ;
        RECT 81.885 42.115 82.055 42.285 ;
        RECT 82.345 42.115 82.515 42.285 ;
        RECT 82.805 42.115 82.975 42.285 ;
        RECT 83.265 42.115 83.435 42.285 ;
        RECT 83.725 42.115 83.895 42.285 ;
        RECT 84.185 42.115 84.355 42.285 ;
        RECT 84.645 42.115 84.815 42.285 ;
        RECT 85.105 42.115 85.275 42.285 ;
        RECT 85.565 42.115 85.735 42.285 ;
        RECT 86.025 42.115 86.195 42.285 ;
        RECT 86.485 42.115 86.655 42.285 ;
        RECT 86.945 42.115 87.115 42.285 ;
        RECT 87.405 42.115 87.575 42.285 ;
        RECT 87.865 42.115 88.035 42.285 ;
        RECT 88.325 42.115 88.495 42.285 ;
        RECT 88.785 42.115 88.955 42.285 ;
        RECT 89.245 42.115 89.415 42.285 ;
        RECT 89.705 42.115 89.875 42.285 ;
        RECT 90.165 42.115 90.335 42.285 ;
        RECT 90.625 42.115 90.795 42.285 ;
        RECT 91.085 42.115 91.255 42.285 ;
        RECT 91.545 42.115 91.715 42.285 ;
        RECT 92.005 42.115 92.175 42.285 ;
        RECT 92.465 42.115 92.635 42.285 ;
        RECT 92.925 42.115 93.095 42.285 ;
        RECT 93.385 42.115 93.555 42.285 ;
        RECT 93.845 42.115 94.015 42.285 ;
        RECT 94.305 42.115 94.475 42.285 ;
        RECT 94.765 42.115 94.935 42.285 ;
        RECT 95.225 42.115 95.395 42.285 ;
        RECT 95.685 42.115 95.855 42.285 ;
        RECT 96.145 42.115 96.315 42.285 ;
        RECT 96.605 42.115 96.775 42.285 ;
        RECT 97.065 42.115 97.235 42.285 ;
        RECT 97.525 42.115 97.695 42.285 ;
        RECT 97.985 42.115 98.155 42.285 ;
        RECT 98.445 42.115 98.615 42.285 ;
        RECT 98.905 42.115 99.075 42.285 ;
        RECT 99.365 42.115 99.535 42.285 ;
        RECT 99.825 42.115 99.995 42.285 ;
        RECT 100.285 42.115 100.455 42.285 ;
        RECT 100.745 42.115 100.915 42.285 ;
        RECT 101.205 42.115 101.375 42.285 ;
        RECT 101.665 42.115 101.835 42.285 ;
        RECT 102.125 42.115 102.295 42.285 ;
        RECT 102.585 42.115 102.755 42.285 ;
        RECT 103.045 42.115 103.215 42.285 ;
        RECT 103.505 42.115 103.675 42.285 ;
        RECT 103.965 42.115 104.135 42.285 ;
        RECT 104.425 42.115 104.595 42.285 ;
        RECT 104.885 42.115 105.055 42.285 ;
        RECT 105.345 42.115 105.515 42.285 ;
        RECT 105.805 42.115 105.975 42.285 ;
        RECT 106.265 42.115 106.435 42.285 ;
        RECT 106.725 42.115 106.895 42.285 ;
        RECT 107.185 42.115 107.355 42.285 ;
        RECT 107.645 42.115 107.815 42.285 ;
        RECT 108.105 42.115 108.275 42.285 ;
        RECT 108.565 42.115 108.735 42.285 ;
        RECT 109.025 42.115 109.195 42.285 ;
        RECT 109.485 42.115 109.655 42.285 ;
        RECT 109.945 42.115 110.115 42.285 ;
        RECT 110.405 42.115 110.575 42.285 ;
        RECT 110.865 42.115 111.035 42.285 ;
        RECT 111.325 42.115 111.495 42.285 ;
        RECT 111.785 42.115 111.955 42.285 ;
        RECT 112.245 42.115 112.415 42.285 ;
        RECT 112.705 42.115 112.875 42.285 ;
        RECT 113.165 42.115 113.335 42.285 ;
        RECT 113.625 42.115 113.795 42.285 ;
        RECT 114.085 42.115 114.255 42.285 ;
        RECT 114.545 42.115 114.715 42.285 ;
        RECT 115.005 42.115 115.175 42.285 ;
        RECT 115.465 42.115 115.635 42.285 ;
        RECT 115.925 42.115 116.095 42.285 ;
        RECT 116.385 42.115 116.555 42.285 ;
        RECT 116.845 42.115 117.015 42.285 ;
        RECT 117.305 42.115 117.475 42.285 ;
        RECT 117.765 42.115 117.935 42.285 ;
        RECT 118.225 42.115 118.395 42.285 ;
        RECT 118.685 42.115 118.855 42.285 ;
        RECT 119.145 42.115 119.315 42.285 ;
        RECT 119.605 42.115 119.775 42.285 ;
        RECT 120.065 42.115 120.235 42.285 ;
        RECT 120.525 42.115 120.695 42.285 ;
        RECT 120.985 42.115 121.155 42.285 ;
        RECT 121.445 42.115 121.615 42.285 ;
        RECT 121.905 42.115 122.075 42.285 ;
        RECT 122.365 42.115 122.535 42.285 ;
        RECT 122.825 42.115 122.995 42.285 ;
        RECT 123.285 42.115 123.455 42.285 ;
        RECT 123.745 42.115 123.915 42.285 ;
        RECT 124.205 42.115 124.375 42.285 ;
        RECT 124.665 42.115 124.835 42.285 ;
        RECT 125.125 42.115 125.295 42.285 ;
        RECT 125.585 42.115 125.755 42.285 ;
        RECT 126.045 42.115 126.215 42.285 ;
        RECT 126.505 42.115 126.675 42.285 ;
        RECT 126.965 42.115 127.135 42.285 ;
        RECT 127.425 42.115 127.595 42.285 ;
        RECT 127.885 42.115 128.055 42.285 ;
        RECT 128.345 42.115 128.515 42.285 ;
        RECT 128.805 42.115 128.975 42.285 ;
        RECT 129.265 42.115 129.435 42.285 ;
        RECT 129.725 42.115 129.895 42.285 ;
        RECT 130.185 42.115 130.355 42.285 ;
        RECT 130.645 42.115 130.815 42.285 ;
        RECT 131.105 42.115 131.275 42.285 ;
        RECT 131.565 42.115 131.735 42.285 ;
        RECT 132.025 42.115 132.195 42.285 ;
        RECT 132.485 42.115 132.655 42.285 ;
        RECT 132.945 42.115 133.115 42.285 ;
        RECT 133.405 42.115 133.575 42.285 ;
        RECT 133.865 42.115 134.035 42.285 ;
        RECT 134.325 42.115 134.495 42.285 ;
        RECT 134.785 42.115 134.955 42.285 ;
        RECT 135.245 42.115 135.415 42.285 ;
        RECT 135.705 42.115 135.875 42.285 ;
        RECT 136.165 42.115 136.335 42.285 ;
        RECT 136.625 42.115 136.795 42.285 ;
        RECT 137.085 42.115 137.255 42.285 ;
        RECT 137.545 42.115 137.715 42.285 ;
        RECT 138.005 42.115 138.175 42.285 ;
        RECT 138.465 42.115 138.635 42.285 ;
        RECT 138.925 42.115 139.095 42.285 ;
        RECT 139.385 42.115 139.555 42.285 ;
        RECT 139.845 42.115 140.015 42.285 ;
        RECT 140.305 42.115 140.475 42.285 ;
        RECT 140.765 42.115 140.935 42.285 ;
        RECT 141.225 42.115 141.395 42.285 ;
        RECT 141.685 42.115 141.855 42.285 ;
        RECT 142.145 42.115 142.315 42.285 ;
        RECT 142.605 42.115 142.775 42.285 ;
        RECT 143.065 42.115 143.235 42.285 ;
        RECT 143.525 42.115 143.695 42.285 ;
        RECT 143.985 42.115 144.155 42.285 ;
        RECT 55.665 36.675 55.835 36.845 ;
        RECT 56.125 36.675 56.295 36.845 ;
        RECT 56.585 36.675 56.755 36.845 ;
        RECT 57.045 36.675 57.215 36.845 ;
        RECT 57.505 36.675 57.675 36.845 ;
        RECT 57.965 36.675 58.135 36.845 ;
        RECT 58.425 36.675 58.595 36.845 ;
        RECT 58.885 36.675 59.055 36.845 ;
        RECT 59.345 36.675 59.515 36.845 ;
        RECT 59.805 36.675 59.975 36.845 ;
        RECT 60.265 36.675 60.435 36.845 ;
        RECT 60.725 36.675 60.895 36.845 ;
        RECT 61.185 36.675 61.355 36.845 ;
        RECT 61.645 36.675 61.815 36.845 ;
        RECT 62.105 36.675 62.275 36.845 ;
        RECT 62.565 36.675 62.735 36.845 ;
        RECT 63.025 36.675 63.195 36.845 ;
        RECT 63.485 36.675 63.655 36.845 ;
        RECT 63.945 36.675 64.115 36.845 ;
        RECT 64.405 36.675 64.575 36.845 ;
        RECT 64.865 36.675 65.035 36.845 ;
        RECT 65.325 36.675 65.495 36.845 ;
        RECT 65.785 36.675 65.955 36.845 ;
        RECT 66.245 36.675 66.415 36.845 ;
        RECT 66.705 36.675 66.875 36.845 ;
        RECT 67.165 36.675 67.335 36.845 ;
        RECT 67.625 36.675 67.795 36.845 ;
        RECT 68.085 36.675 68.255 36.845 ;
        RECT 68.545 36.675 68.715 36.845 ;
        RECT 69.005 36.675 69.175 36.845 ;
        RECT 69.465 36.675 69.635 36.845 ;
        RECT 69.925 36.675 70.095 36.845 ;
        RECT 70.385 36.675 70.555 36.845 ;
        RECT 70.845 36.675 71.015 36.845 ;
        RECT 71.305 36.675 71.475 36.845 ;
        RECT 71.765 36.675 71.935 36.845 ;
        RECT 72.225 36.675 72.395 36.845 ;
        RECT 72.685 36.675 72.855 36.845 ;
        RECT 73.145 36.675 73.315 36.845 ;
        RECT 73.605 36.675 73.775 36.845 ;
        RECT 74.065 36.675 74.235 36.845 ;
        RECT 74.525 36.675 74.695 36.845 ;
        RECT 74.985 36.675 75.155 36.845 ;
        RECT 75.445 36.675 75.615 36.845 ;
        RECT 75.905 36.675 76.075 36.845 ;
        RECT 76.365 36.675 76.535 36.845 ;
        RECT 76.825 36.675 76.995 36.845 ;
        RECT 77.285 36.675 77.455 36.845 ;
        RECT 77.745 36.675 77.915 36.845 ;
        RECT 78.205 36.675 78.375 36.845 ;
        RECT 78.665 36.675 78.835 36.845 ;
        RECT 79.125 36.675 79.295 36.845 ;
        RECT 79.585 36.675 79.755 36.845 ;
        RECT 80.045 36.675 80.215 36.845 ;
        RECT 80.505 36.675 80.675 36.845 ;
        RECT 80.965 36.675 81.135 36.845 ;
        RECT 81.425 36.675 81.595 36.845 ;
        RECT 81.885 36.675 82.055 36.845 ;
        RECT 82.345 36.675 82.515 36.845 ;
        RECT 82.805 36.675 82.975 36.845 ;
        RECT 83.265 36.675 83.435 36.845 ;
        RECT 83.725 36.675 83.895 36.845 ;
        RECT 84.185 36.675 84.355 36.845 ;
        RECT 84.645 36.675 84.815 36.845 ;
        RECT 85.105 36.675 85.275 36.845 ;
        RECT 85.565 36.675 85.735 36.845 ;
        RECT 86.025 36.675 86.195 36.845 ;
        RECT 86.485 36.675 86.655 36.845 ;
        RECT 86.945 36.675 87.115 36.845 ;
        RECT 87.405 36.675 87.575 36.845 ;
        RECT 87.865 36.675 88.035 36.845 ;
        RECT 88.325 36.675 88.495 36.845 ;
        RECT 88.785 36.675 88.955 36.845 ;
        RECT 89.245 36.675 89.415 36.845 ;
        RECT 89.705 36.675 89.875 36.845 ;
        RECT 90.165 36.675 90.335 36.845 ;
        RECT 90.625 36.675 90.795 36.845 ;
        RECT 91.085 36.675 91.255 36.845 ;
        RECT 91.545 36.675 91.715 36.845 ;
        RECT 92.005 36.675 92.175 36.845 ;
        RECT 92.465 36.675 92.635 36.845 ;
        RECT 92.925 36.675 93.095 36.845 ;
        RECT 93.385 36.675 93.555 36.845 ;
        RECT 93.845 36.675 94.015 36.845 ;
        RECT 94.305 36.675 94.475 36.845 ;
        RECT 94.765 36.675 94.935 36.845 ;
        RECT 95.225 36.675 95.395 36.845 ;
        RECT 95.685 36.675 95.855 36.845 ;
        RECT 96.145 36.675 96.315 36.845 ;
        RECT 96.605 36.675 96.775 36.845 ;
        RECT 97.065 36.675 97.235 36.845 ;
        RECT 97.525 36.675 97.695 36.845 ;
        RECT 97.985 36.675 98.155 36.845 ;
        RECT 98.445 36.675 98.615 36.845 ;
        RECT 98.905 36.675 99.075 36.845 ;
        RECT 99.365 36.675 99.535 36.845 ;
        RECT 99.825 36.675 99.995 36.845 ;
        RECT 100.285 36.675 100.455 36.845 ;
        RECT 100.745 36.675 100.915 36.845 ;
        RECT 101.205 36.675 101.375 36.845 ;
        RECT 101.665 36.675 101.835 36.845 ;
        RECT 102.125 36.675 102.295 36.845 ;
        RECT 102.585 36.675 102.755 36.845 ;
        RECT 103.045 36.675 103.215 36.845 ;
        RECT 103.505 36.675 103.675 36.845 ;
        RECT 103.965 36.675 104.135 36.845 ;
        RECT 104.425 36.675 104.595 36.845 ;
        RECT 104.885 36.675 105.055 36.845 ;
        RECT 105.345 36.675 105.515 36.845 ;
        RECT 105.805 36.675 105.975 36.845 ;
        RECT 106.265 36.675 106.435 36.845 ;
        RECT 106.725 36.675 106.895 36.845 ;
        RECT 107.185 36.675 107.355 36.845 ;
        RECT 107.645 36.675 107.815 36.845 ;
        RECT 108.105 36.675 108.275 36.845 ;
        RECT 108.565 36.675 108.735 36.845 ;
        RECT 109.025 36.675 109.195 36.845 ;
        RECT 109.485 36.675 109.655 36.845 ;
        RECT 109.945 36.675 110.115 36.845 ;
        RECT 110.405 36.675 110.575 36.845 ;
        RECT 110.865 36.675 111.035 36.845 ;
        RECT 111.325 36.675 111.495 36.845 ;
        RECT 111.785 36.675 111.955 36.845 ;
        RECT 112.245 36.675 112.415 36.845 ;
        RECT 112.705 36.675 112.875 36.845 ;
        RECT 113.165 36.675 113.335 36.845 ;
        RECT 113.625 36.675 113.795 36.845 ;
        RECT 114.085 36.675 114.255 36.845 ;
        RECT 114.545 36.675 114.715 36.845 ;
        RECT 115.005 36.675 115.175 36.845 ;
        RECT 115.465 36.675 115.635 36.845 ;
        RECT 115.925 36.675 116.095 36.845 ;
        RECT 116.385 36.675 116.555 36.845 ;
        RECT 116.845 36.675 117.015 36.845 ;
        RECT 117.305 36.675 117.475 36.845 ;
        RECT 117.765 36.675 117.935 36.845 ;
        RECT 118.225 36.675 118.395 36.845 ;
        RECT 118.685 36.675 118.855 36.845 ;
        RECT 119.145 36.675 119.315 36.845 ;
        RECT 119.605 36.675 119.775 36.845 ;
        RECT 120.065 36.675 120.235 36.845 ;
        RECT 120.525 36.675 120.695 36.845 ;
        RECT 120.985 36.675 121.155 36.845 ;
        RECT 121.445 36.675 121.615 36.845 ;
        RECT 121.905 36.675 122.075 36.845 ;
        RECT 122.365 36.675 122.535 36.845 ;
        RECT 122.825 36.675 122.995 36.845 ;
        RECT 123.285 36.675 123.455 36.845 ;
        RECT 123.745 36.675 123.915 36.845 ;
        RECT 124.205 36.675 124.375 36.845 ;
        RECT 124.665 36.675 124.835 36.845 ;
        RECT 125.125 36.675 125.295 36.845 ;
        RECT 125.585 36.675 125.755 36.845 ;
        RECT 126.045 36.675 126.215 36.845 ;
        RECT 126.505 36.675 126.675 36.845 ;
        RECT 126.965 36.675 127.135 36.845 ;
        RECT 127.425 36.675 127.595 36.845 ;
        RECT 127.885 36.675 128.055 36.845 ;
        RECT 128.345 36.675 128.515 36.845 ;
        RECT 128.805 36.675 128.975 36.845 ;
        RECT 129.265 36.675 129.435 36.845 ;
        RECT 129.725 36.675 129.895 36.845 ;
        RECT 130.185 36.675 130.355 36.845 ;
        RECT 130.645 36.675 130.815 36.845 ;
        RECT 131.105 36.675 131.275 36.845 ;
        RECT 131.565 36.675 131.735 36.845 ;
        RECT 132.025 36.675 132.195 36.845 ;
        RECT 132.485 36.675 132.655 36.845 ;
        RECT 132.945 36.675 133.115 36.845 ;
        RECT 133.405 36.675 133.575 36.845 ;
        RECT 133.865 36.675 134.035 36.845 ;
        RECT 134.325 36.675 134.495 36.845 ;
        RECT 134.785 36.675 134.955 36.845 ;
        RECT 135.245 36.675 135.415 36.845 ;
        RECT 135.705 36.675 135.875 36.845 ;
        RECT 136.165 36.675 136.335 36.845 ;
        RECT 136.625 36.675 136.795 36.845 ;
        RECT 137.085 36.675 137.255 36.845 ;
        RECT 137.545 36.675 137.715 36.845 ;
        RECT 138.005 36.675 138.175 36.845 ;
        RECT 138.465 36.675 138.635 36.845 ;
        RECT 138.925 36.675 139.095 36.845 ;
        RECT 139.385 36.675 139.555 36.845 ;
        RECT 139.845 36.675 140.015 36.845 ;
        RECT 140.305 36.675 140.475 36.845 ;
        RECT 140.765 36.675 140.935 36.845 ;
        RECT 141.225 36.675 141.395 36.845 ;
        RECT 141.685 36.675 141.855 36.845 ;
        RECT 142.145 36.675 142.315 36.845 ;
        RECT 142.605 36.675 142.775 36.845 ;
        RECT 143.065 36.675 143.235 36.845 ;
        RECT 143.525 36.675 143.695 36.845 ;
        RECT 143.985 36.675 144.155 36.845 ;
        RECT 55.665 31.235 55.835 31.405 ;
        RECT 56.125 31.235 56.295 31.405 ;
        RECT 56.585 31.235 56.755 31.405 ;
        RECT 57.045 31.235 57.215 31.405 ;
        RECT 57.505 31.235 57.675 31.405 ;
        RECT 57.965 31.235 58.135 31.405 ;
        RECT 58.425 31.235 58.595 31.405 ;
        RECT 58.885 31.235 59.055 31.405 ;
        RECT 59.345 31.235 59.515 31.405 ;
        RECT 59.805 31.235 59.975 31.405 ;
        RECT 60.265 31.235 60.435 31.405 ;
        RECT 60.725 31.235 60.895 31.405 ;
        RECT 61.185 31.235 61.355 31.405 ;
        RECT 61.645 31.235 61.815 31.405 ;
        RECT 62.105 31.235 62.275 31.405 ;
        RECT 62.565 31.235 62.735 31.405 ;
        RECT 63.025 31.235 63.195 31.405 ;
        RECT 63.485 31.235 63.655 31.405 ;
        RECT 63.945 31.235 64.115 31.405 ;
        RECT 64.405 31.235 64.575 31.405 ;
        RECT 64.865 31.235 65.035 31.405 ;
        RECT 65.325 31.235 65.495 31.405 ;
        RECT 65.785 31.235 65.955 31.405 ;
        RECT 66.245 31.235 66.415 31.405 ;
        RECT 66.705 31.235 66.875 31.405 ;
        RECT 67.165 31.235 67.335 31.405 ;
        RECT 67.625 31.235 67.795 31.405 ;
        RECT 68.085 31.235 68.255 31.405 ;
        RECT 68.545 31.235 68.715 31.405 ;
        RECT 69.005 31.235 69.175 31.405 ;
        RECT 69.465 31.235 69.635 31.405 ;
        RECT 69.925 31.235 70.095 31.405 ;
        RECT 70.385 31.235 70.555 31.405 ;
        RECT 70.845 31.235 71.015 31.405 ;
        RECT 71.305 31.235 71.475 31.405 ;
        RECT 71.765 31.235 71.935 31.405 ;
        RECT 72.225 31.235 72.395 31.405 ;
        RECT 72.685 31.235 72.855 31.405 ;
        RECT 73.145 31.235 73.315 31.405 ;
        RECT 73.605 31.235 73.775 31.405 ;
        RECT 74.065 31.235 74.235 31.405 ;
        RECT 74.525 31.235 74.695 31.405 ;
        RECT 74.985 31.235 75.155 31.405 ;
        RECT 75.445 31.235 75.615 31.405 ;
        RECT 75.905 31.235 76.075 31.405 ;
        RECT 76.365 31.235 76.535 31.405 ;
        RECT 76.825 31.235 76.995 31.405 ;
        RECT 77.285 31.235 77.455 31.405 ;
        RECT 77.745 31.235 77.915 31.405 ;
        RECT 78.205 31.235 78.375 31.405 ;
        RECT 78.665 31.235 78.835 31.405 ;
        RECT 79.125 31.235 79.295 31.405 ;
        RECT 79.585 31.235 79.755 31.405 ;
        RECT 80.045 31.235 80.215 31.405 ;
        RECT 80.505 31.235 80.675 31.405 ;
        RECT 80.965 31.235 81.135 31.405 ;
        RECT 81.425 31.235 81.595 31.405 ;
        RECT 81.885 31.235 82.055 31.405 ;
        RECT 82.345 31.235 82.515 31.405 ;
        RECT 82.805 31.235 82.975 31.405 ;
        RECT 83.265 31.235 83.435 31.405 ;
        RECT 83.725 31.235 83.895 31.405 ;
        RECT 84.185 31.235 84.355 31.405 ;
        RECT 84.645 31.235 84.815 31.405 ;
        RECT 85.105 31.235 85.275 31.405 ;
        RECT 85.565 31.235 85.735 31.405 ;
        RECT 86.025 31.235 86.195 31.405 ;
        RECT 86.485 31.235 86.655 31.405 ;
        RECT 86.945 31.235 87.115 31.405 ;
        RECT 87.405 31.235 87.575 31.405 ;
        RECT 87.865 31.235 88.035 31.405 ;
        RECT 88.325 31.235 88.495 31.405 ;
        RECT 88.785 31.235 88.955 31.405 ;
        RECT 89.245 31.235 89.415 31.405 ;
        RECT 89.705 31.235 89.875 31.405 ;
        RECT 90.165 31.235 90.335 31.405 ;
        RECT 90.625 31.235 90.795 31.405 ;
        RECT 91.085 31.235 91.255 31.405 ;
        RECT 91.545 31.235 91.715 31.405 ;
        RECT 92.005 31.235 92.175 31.405 ;
        RECT 92.465 31.235 92.635 31.405 ;
        RECT 92.925 31.235 93.095 31.405 ;
        RECT 93.385 31.235 93.555 31.405 ;
        RECT 93.845 31.235 94.015 31.405 ;
        RECT 94.305 31.235 94.475 31.405 ;
        RECT 94.765 31.235 94.935 31.405 ;
        RECT 95.225 31.235 95.395 31.405 ;
        RECT 95.685 31.235 95.855 31.405 ;
        RECT 96.145 31.235 96.315 31.405 ;
        RECT 96.605 31.235 96.775 31.405 ;
        RECT 97.065 31.235 97.235 31.405 ;
        RECT 97.525 31.235 97.695 31.405 ;
        RECT 97.985 31.235 98.155 31.405 ;
        RECT 98.445 31.235 98.615 31.405 ;
        RECT 98.905 31.235 99.075 31.405 ;
        RECT 99.365 31.235 99.535 31.405 ;
        RECT 99.825 31.235 99.995 31.405 ;
        RECT 100.285 31.235 100.455 31.405 ;
        RECT 100.745 31.235 100.915 31.405 ;
        RECT 101.205 31.235 101.375 31.405 ;
        RECT 101.665 31.235 101.835 31.405 ;
        RECT 102.125 31.235 102.295 31.405 ;
        RECT 102.585 31.235 102.755 31.405 ;
        RECT 103.045 31.235 103.215 31.405 ;
        RECT 103.505 31.235 103.675 31.405 ;
        RECT 103.965 31.235 104.135 31.405 ;
        RECT 104.425 31.235 104.595 31.405 ;
        RECT 104.885 31.235 105.055 31.405 ;
        RECT 105.345 31.235 105.515 31.405 ;
        RECT 105.805 31.235 105.975 31.405 ;
        RECT 106.265 31.235 106.435 31.405 ;
        RECT 106.725 31.235 106.895 31.405 ;
        RECT 107.185 31.235 107.355 31.405 ;
        RECT 107.645 31.235 107.815 31.405 ;
        RECT 108.105 31.235 108.275 31.405 ;
        RECT 108.565 31.235 108.735 31.405 ;
        RECT 109.025 31.235 109.195 31.405 ;
        RECT 109.485 31.235 109.655 31.405 ;
        RECT 109.945 31.235 110.115 31.405 ;
        RECT 110.405 31.235 110.575 31.405 ;
        RECT 110.865 31.235 111.035 31.405 ;
        RECT 111.325 31.235 111.495 31.405 ;
        RECT 111.785 31.235 111.955 31.405 ;
        RECT 112.245 31.235 112.415 31.405 ;
        RECT 112.705 31.235 112.875 31.405 ;
        RECT 113.165 31.235 113.335 31.405 ;
        RECT 113.625 31.235 113.795 31.405 ;
        RECT 114.085 31.235 114.255 31.405 ;
        RECT 114.545 31.235 114.715 31.405 ;
        RECT 115.005 31.235 115.175 31.405 ;
        RECT 115.465 31.235 115.635 31.405 ;
        RECT 115.925 31.235 116.095 31.405 ;
        RECT 116.385 31.235 116.555 31.405 ;
        RECT 116.845 31.235 117.015 31.405 ;
        RECT 117.305 31.235 117.475 31.405 ;
        RECT 117.765 31.235 117.935 31.405 ;
        RECT 118.225 31.235 118.395 31.405 ;
        RECT 118.685 31.235 118.855 31.405 ;
        RECT 119.145 31.235 119.315 31.405 ;
        RECT 119.605 31.235 119.775 31.405 ;
        RECT 120.065 31.235 120.235 31.405 ;
        RECT 120.525 31.235 120.695 31.405 ;
        RECT 120.985 31.235 121.155 31.405 ;
        RECT 121.445 31.235 121.615 31.405 ;
        RECT 121.905 31.235 122.075 31.405 ;
        RECT 122.365 31.235 122.535 31.405 ;
        RECT 122.825 31.235 122.995 31.405 ;
        RECT 123.285 31.235 123.455 31.405 ;
        RECT 123.745 31.235 123.915 31.405 ;
        RECT 124.205 31.235 124.375 31.405 ;
        RECT 124.665 31.235 124.835 31.405 ;
        RECT 125.125 31.235 125.295 31.405 ;
        RECT 125.585 31.235 125.755 31.405 ;
        RECT 126.045 31.235 126.215 31.405 ;
        RECT 126.505 31.235 126.675 31.405 ;
        RECT 126.965 31.235 127.135 31.405 ;
        RECT 127.425 31.235 127.595 31.405 ;
        RECT 127.885 31.235 128.055 31.405 ;
        RECT 128.345 31.235 128.515 31.405 ;
        RECT 128.805 31.235 128.975 31.405 ;
        RECT 129.265 31.235 129.435 31.405 ;
        RECT 129.725 31.235 129.895 31.405 ;
        RECT 130.185 31.235 130.355 31.405 ;
        RECT 130.645 31.235 130.815 31.405 ;
        RECT 131.105 31.235 131.275 31.405 ;
        RECT 131.565 31.235 131.735 31.405 ;
        RECT 132.025 31.235 132.195 31.405 ;
        RECT 132.485 31.235 132.655 31.405 ;
        RECT 132.945 31.235 133.115 31.405 ;
        RECT 133.405 31.235 133.575 31.405 ;
        RECT 133.865 31.235 134.035 31.405 ;
        RECT 134.325 31.235 134.495 31.405 ;
        RECT 134.785 31.235 134.955 31.405 ;
        RECT 135.245 31.235 135.415 31.405 ;
        RECT 135.705 31.235 135.875 31.405 ;
        RECT 136.165 31.235 136.335 31.405 ;
        RECT 136.625 31.235 136.795 31.405 ;
        RECT 137.085 31.235 137.255 31.405 ;
        RECT 137.545 31.235 137.715 31.405 ;
        RECT 138.005 31.235 138.175 31.405 ;
        RECT 138.465 31.235 138.635 31.405 ;
        RECT 138.925 31.235 139.095 31.405 ;
        RECT 139.385 31.235 139.555 31.405 ;
        RECT 139.845 31.235 140.015 31.405 ;
        RECT 140.305 31.235 140.475 31.405 ;
        RECT 140.765 31.235 140.935 31.405 ;
        RECT 141.225 31.235 141.395 31.405 ;
        RECT 141.685 31.235 141.855 31.405 ;
        RECT 142.145 31.235 142.315 31.405 ;
        RECT 142.605 31.235 142.775 31.405 ;
        RECT 143.065 31.235 143.235 31.405 ;
        RECT 143.525 31.235 143.695 31.405 ;
        RECT 143.985 31.235 144.155 31.405 ;
        RECT 55.665 25.795 55.835 25.965 ;
        RECT 56.125 25.795 56.295 25.965 ;
        RECT 56.585 25.795 56.755 25.965 ;
        RECT 57.045 25.795 57.215 25.965 ;
        RECT 57.505 25.795 57.675 25.965 ;
        RECT 57.965 25.795 58.135 25.965 ;
        RECT 58.425 25.795 58.595 25.965 ;
        RECT 58.885 25.795 59.055 25.965 ;
        RECT 59.345 25.795 59.515 25.965 ;
        RECT 59.805 25.795 59.975 25.965 ;
        RECT 60.265 25.795 60.435 25.965 ;
        RECT 60.725 25.795 60.895 25.965 ;
        RECT 61.185 25.795 61.355 25.965 ;
        RECT 61.645 25.795 61.815 25.965 ;
        RECT 62.105 25.795 62.275 25.965 ;
        RECT 62.565 25.795 62.735 25.965 ;
        RECT 63.025 25.795 63.195 25.965 ;
        RECT 63.485 25.795 63.655 25.965 ;
        RECT 63.945 25.795 64.115 25.965 ;
        RECT 64.405 25.795 64.575 25.965 ;
        RECT 64.865 25.795 65.035 25.965 ;
        RECT 65.325 25.795 65.495 25.965 ;
        RECT 65.785 25.795 65.955 25.965 ;
        RECT 66.245 25.795 66.415 25.965 ;
        RECT 66.705 25.795 66.875 25.965 ;
        RECT 67.165 25.795 67.335 25.965 ;
        RECT 67.625 25.795 67.795 25.965 ;
        RECT 68.085 25.795 68.255 25.965 ;
        RECT 68.545 25.795 68.715 25.965 ;
        RECT 69.005 25.795 69.175 25.965 ;
        RECT 69.465 25.795 69.635 25.965 ;
        RECT 69.925 25.795 70.095 25.965 ;
        RECT 70.385 25.795 70.555 25.965 ;
        RECT 70.845 25.795 71.015 25.965 ;
        RECT 71.305 25.795 71.475 25.965 ;
        RECT 71.765 25.795 71.935 25.965 ;
        RECT 72.225 25.795 72.395 25.965 ;
        RECT 72.685 25.795 72.855 25.965 ;
        RECT 73.145 25.795 73.315 25.965 ;
        RECT 73.605 25.795 73.775 25.965 ;
        RECT 74.065 25.795 74.235 25.965 ;
        RECT 74.525 25.795 74.695 25.965 ;
        RECT 74.985 25.795 75.155 25.965 ;
        RECT 75.445 25.795 75.615 25.965 ;
        RECT 75.905 25.795 76.075 25.965 ;
        RECT 76.365 25.795 76.535 25.965 ;
        RECT 76.825 25.795 76.995 25.965 ;
        RECT 77.285 25.795 77.455 25.965 ;
        RECT 77.745 25.795 77.915 25.965 ;
        RECT 78.205 25.795 78.375 25.965 ;
        RECT 78.665 25.795 78.835 25.965 ;
        RECT 79.125 25.795 79.295 25.965 ;
        RECT 79.585 25.795 79.755 25.965 ;
        RECT 80.045 25.795 80.215 25.965 ;
        RECT 80.505 25.795 80.675 25.965 ;
        RECT 80.965 25.795 81.135 25.965 ;
        RECT 81.425 25.795 81.595 25.965 ;
        RECT 81.885 25.795 82.055 25.965 ;
        RECT 82.345 25.795 82.515 25.965 ;
        RECT 82.805 25.795 82.975 25.965 ;
        RECT 83.265 25.795 83.435 25.965 ;
        RECT 83.725 25.795 83.895 25.965 ;
        RECT 84.185 25.795 84.355 25.965 ;
        RECT 84.645 25.795 84.815 25.965 ;
        RECT 85.105 25.795 85.275 25.965 ;
        RECT 85.565 25.795 85.735 25.965 ;
        RECT 86.025 25.795 86.195 25.965 ;
        RECT 86.485 25.795 86.655 25.965 ;
        RECT 86.945 25.795 87.115 25.965 ;
        RECT 87.405 25.795 87.575 25.965 ;
        RECT 87.865 25.795 88.035 25.965 ;
        RECT 88.325 25.795 88.495 25.965 ;
        RECT 88.785 25.795 88.955 25.965 ;
        RECT 89.245 25.795 89.415 25.965 ;
        RECT 89.705 25.795 89.875 25.965 ;
        RECT 90.165 25.795 90.335 25.965 ;
        RECT 90.625 25.795 90.795 25.965 ;
        RECT 91.085 25.795 91.255 25.965 ;
        RECT 91.545 25.795 91.715 25.965 ;
        RECT 92.005 25.795 92.175 25.965 ;
        RECT 92.465 25.795 92.635 25.965 ;
        RECT 92.925 25.795 93.095 25.965 ;
        RECT 93.385 25.795 93.555 25.965 ;
        RECT 93.845 25.795 94.015 25.965 ;
        RECT 94.305 25.795 94.475 25.965 ;
        RECT 94.765 25.795 94.935 25.965 ;
        RECT 95.225 25.795 95.395 25.965 ;
        RECT 95.685 25.795 95.855 25.965 ;
        RECT 96.145 25.795 96.315 25.965 ;
        RECT 96.605 25.795 96.775 25.965 ;
        RECT 97.065 25.795 97.235 25.965 ;
        RECT 97.525 25.795 97.695 25.965 ;
        RECT 97.985 25.795 98.155 25.965 ;
        RECT 98.445 25.795 98.615 25.965 ;
        RECT 98.905 25.795 99.075 25.965 ;
        RECT 99.365 25.795 99.535 25.965 ;
        RECT 99.825 25.795 99.995 25.965 ;
        RECT 100.285 25.795 100.455 25.965 ;
        RECT 100.745 25.795 100.915 25.965 ;
        RECT 101.205 25.795 101.375 25.965 ;
        RECT 101.665 25.795 101.835 25.965 ;
        RECT 102.125 25.795 102.295 25.965 ;
        RECT 102.585 25.795 102.755 25.965 ;
        RECT 103.045 25.795 103.215 25.965 ;
        RECT 103.505 25.795 103.675 25.965 ;
        RECT 103.965 25.795 104.135 25.965 ;
        RECT 104.425 25.795 104.595 25.965 ;
        RECT 104.885 25.795 105.055 25.965 ;
        RECT 105.345 25.795 105.515 25.965 ;
        RECT 105.805 25.795 105.975 25.965 ;
        RECT 106.265 25.795 106.435 25.965 ;
        RECT 106.725 25.795 106.895 25.965 ;
        RECT 107.185 25.795 107.355 25.965 ;
        RECT 107.645 25.795 107.815 25.965 ;
        RECT 108.105 25.795 108.275 25.965 ;
        RECT 108.565 25.795 108.735 25.965 ;
        RECT 109.025 25.795 109.195 25.965 ;
        RECT 109.485 25.795 109.655 25.965 ;
        RECT 109.945 25.795 110.115 25.965 ;
        RECT 110.405 25.795 110.575 25.965 ;
        RECT 110.865 25.795 111.035 25.965 ;
        RECT 111.325 25.795 111.495 25.965 ;
        RECT 111.785 25.795 111.955 25.965 ;
        RECT 112.245 25.795 112.415 25.965 ;
        RECT 112.705 25.795 112.875 25.965 ;
        RECT 113.165 25.795 113.335 25.965 ;
        RECT 113.625 25.795 113.795 25.965 ;
        RECT 114.085 25.795 114.255 25.965 ;
        RECT 114.545 25.795 114.715 25.965 ;
        RECT 115.005 25.795 115.175 25.965 ;
        RECT 115.465 25.795 115.635 25.965 ;
        RECT 115.925 25.795 116.095 25.965 ;
        RECT 116.385 25.795 116.555 25.965 ;
        RECT 116.845 25.795 117.015 25.965 ;
        RECT 117.305 25.795 117.475 25.965 ;
        RECT 117.765 25.795 117.935 25.965 ;
        RECT 118.225 25.795 118.395 25.965 ;
        RECT 118.685 25.795 118.855 25.965 ;
        RECT 119.145 25.795 119.315 25.965 ;
        RECT 119.605 25.795 119.775 25.965 ;
        RECT 120.065 25.795 120.235 25.965 ;
        RECT 120.525 25.795 120.695 25.965 ;
        RECT 120.985 25.795 121.155 25.965 ;
        RECT 121.445 25.795 121.615 25.965 ;
        RECT 121.905 25.795 122.075 25.965 ;
        RECT 122.365 25.795 122.535 25.965 ;
        RECT 122.825 25.795 122.995 25.965 ;
        RECT 123.285 25.795 123.455 25.965 ;
        RECT 123.745 25.795 123.915 25.965 ;
        RECT 124.205 25.795 124.375 25.965 ;
        RECT 124.665 25.795 124.835 25.965 ;
        RECT 125.125 25.795 125.295 25.965 ;
        RECT 125.585 25.795 125.755 25.965 ;
        RECT 126.045 25.795 126.215 25.965 ;
        RECT 126.505 25.795 126.675 25.965 ;
        RECT 126.965 25.795 127.135 25.965 ;
        RECT 127.425 25.795 127.595 25.965 ;
        RECT 127.885 25.795 128.055 25.965 ;
        RECT 128.345 25.795 128.515 25.965 ;
        RECT 128.805 25.795 128.975 25.965 ;
        RECT 129.265 25.795 129.435 25.965 ;
        RECT 129.725 25.795 129.895 25.965 ;
        RECT 130.185 25.795 130.355 25.965 ;
        RECT 130.645 25.795 130.815 25.965 ;
        RECT 131.105 25.795 131.275 25.965 ;
        RECT 131.565 25.795 131.735 25.965 ;
        RECT 132.025 25.795 132.195 25.965 ;
        RECT 132.485 25.795 132.655 25.965 ;
        RECT 132.945 25.795 133.115 25.965 ;
        RECT 133.405 25.795 133.575 25.965 ;
        RECT 133.865 25.795 134.035 25.965 ;
        RECT 134.325 25.795 134.495 25.965 ;
        RECT 134.785 25.795 134.955 25.965 ;
        RECT 135.245 25.795 135.415 25.965 ;
        RECT 135.705 25.795 135.875 25.965 ;
        RECT 136.165 25.795 136.335 25.965 ;
        RECT 136.625 25.795 136.795 25.965 ;
        RECT 137.085 25.795 137.255 25.965 ;
        RECT 137.545 25.795 137.715 25.965 ;
        RECT 138.005 25.795 138.175 25.965 ;
        RECT 138.465 25.795 138.635 25.965 ;
        RECT 138.925 25.795 139.095 25.965 ;
        RECT 139.385 25.795 139.555 25.965 ;
        RECT 139.845 25.795 140.015 25.965 ;
        RECT 140.305 25.795 140.475 25.965 ;
        RECT 140.765 25.795 140.935 25.965 ;
        RECT 141.225 25.795 141.395 25.965 ;
        RECT 141.685 25.795 141.855 25.965 ;
        RECT 142.145 25.795 142.315 25.965 ;
        RECT 142.605 25.795 142.775 25.965 ;
        RECT 143.065 25.795 143.235 25.965 ;
        RECT 143.525 25.795 143.695 25.965 ;
        RECT 143.985 25.795 144.155 25.965 ;
      LAYER met1 ;
        RECT 55.520 101.800 145.095 102.280 ;
        RECT 55.520 96.360 145.095 96.840 ;
        RECT 55.520 90.920 145.095 91.400 ;
        RECT 55.520 85.480 145.095 85.960 ;
        RECT 55.520 80.040 145.095 80.520 ;
        RECT 55.520 74.600 145.095 75.080 ;
        RECT 55.520 69.160 145.095 69.640 ;
        RECT 55.520 63.720 145.095 64.200 ;
        RECT 55.520 58.280 145.095 58.760 ;
        RECT 55.520 52.840 145.095 53.320 ;
        RECT 55.520 47.400 145.095 47.880 ;
        RECT 55.520 41.960 145.095 42.440 ;
        RECT 55.520 36.520 145.095 37.000 ;
        RECT 55.520 31.080 145.095 31.560 ;
        RECT 55.520 25.640 145.095 26.120 ;
      LAYER via ;
        RECT 76.940 101.910 77.200 102.170 ;
        RECT 77.260 101.910 77.520 102.170 ;
        RECT 77.580 101.910 77.840 102.170 ;
        RECT 77.900 101.910 78.160 102.170 ;
        RECT 78.220 101.910 78.480 102.170 ;
        RECT 99.135 101.910 99.395 102.170 ;
        RECT 99.455 101.910 99.715 102.170 ;
        RECT 99.775 101.910 100.035 102.170 ;
        RECT 100.095 101.910 100.355 102.170 ;
        RECT 100.415 101.910 100.675 102.170 ;
        RECT 121.330 101.910 121.590 102.170 ;
        RECT 121.650 101.910 121.910 102.170 ;
        RECT 121.970 101.910 122.230 102.170 ;
        RECT 122.290 101.910 122.550 102.170 ;
        RECT 122.610 101.910 122.870 102.170 ;
        RECT 143.525 101.910 143.785 102.170 ;
        RECT 143.845 101.910 144.105 102.170 ;
        RECT 144.165 101.910 144.425 102.170 ;
        RECT 144.485 101.910 144.745 102.170 ;
        RECT 144.805 101.910 145.065 102.170 ;
        RECT 76.940 96.470 77.200 96.730 ;
        RECT 77.260 96.470 77.520 96.730 ;
        RECT 77.580 96.470 77.840 96.730 ;
        RECT 77.900 96.470 78.160 96.730 ;
        RECT 78.220 96.470 78.480 96.730 ;
        RECT 99.135 96.470 99.395 96.730 ;
        RECT 99.455 96.470 99.715 96.730 ;
        RECT 99.775 96.470 100.035 96.730 ;
        RECT 100.095 96.470 100.355 96.730 ;
        RECT 100.415 96.470 100.675 96.730 ;
        RECT 121.330 96.470 121.590 96.730 ;
        RECT 121.650 96.470 121.910 96.730 ;
        RECT 121.970 96.470 122.230 96.730 ;
        RECT 122.290 96.470 122.550 96.730 ;
        RECT 122.610 96.470 122.870 96.730 ;
        RECT 143.525 96.470 143.785 96.730 ;
        RECT 143.845 96.470 144.105 96.730 ;
        RECT 144.165 96.470 144.425 96.730 ;
        RECT 144.485 96.470 144.745 96.730 ;
        RECT 144.805 96.470 145.065 96.730 ;
        RECT 76.940 91.030 77.200 91.290 ;
        RECT 77.260 91.030 77.520 91.290 ;
        RECT 77.580 91.030 77.840 91.290 ;
        RECT 77.900 91.030 78.160 91.290 ;
        RECT 78.220 91.030 78.480 91.290 ;
        RECT 99.135 91.030 99.395 91.290 ;
        RECT 99.455 91.030 99.715 91.290 ;
        RECT 99.775 91.030 100.035 91.290 ;
        RECT 100.095 91.030 100.355 91.290 ;
        RECT 100.415 91.030 100.675 91.290 ;
        RECT 121.330 91.030 121.590 91.290 ;
        RECT 121.650 91.030 121.910 91.290 ;
        RECT 121.970 91.030 122.230 91.290 ;
        RECT 122.290 91.030 122.550 91.290 ;
        RECT 122.610 91.030 122.870 91.290 ;
        RECT 143.525 91.030 143.785 91.290 ;
        RECT 143.845 91.030 144.105 91.290 ;
        RECT 144.165 91.030 144.425 91.290 ;
        RECT 144.485 91.030 144.745 91.290 ;
        RECT 144.805 91.030 145.065 91.290 ;
        RECT 76.940 85.590 77.200 85.850 ;
        RECT 77.260 85.590 77.520 85.850 ;
        RECT 77.580 85.590 77.840 85.850 ;
        RECT 77.900 85.590 78.160 85.850 ;
        RECT 78.220 85.590 78.480 85.850 ;
        RECT 99.135 85.590 99.395 85.850 ;
        RECT 99.455 85.590 99.715 85.850 ;
        RECT 99.775 85.590 100.035 85.850 ;
        RECT 100.095 85.590 100.355 85.850 ;
        RECT 100.415 85.590 100.675 85.850 ;
        RECT 121.330 85.590 121.590 85.850 ;
        RECT 121.650 85.590 121.910 85.850 ;
        RECT 121.970 85.590 122.230 85.850 ;
        RECT 122.290 85.590 122.550 85.850 ;
        RECT 122.610 85.590 122.870 85.850 ;
        RECT 143.525 85.590 143.785 85.850 ;
        RECT 143.845 85.590 144.105 85.850 ;
        RECT 144.165 85.590 144.425 85.850 ;
        RECT 144.485 85.590 144.745 85.850 ;
        RECT 144.805 85.590 145.065 85.850 ;
        RECT 76.940 80.150 77.200 80.410 ;
        RECT 77.260 80.150 77.520 80.410 ;
        RECT 77.580 80.150 77.840 80.410 ;
        RECT 77.900 80.150 78.160 80.410 ;
        RECT 78.220 80.150 78.480 80.410 ;
        RECT 99.135 80.150 99.395 80.410 ;
        RECT 99.455 80.150 99.715 80.410 ;
        RECT 99.775 80.150 100.035 80.410 ;
        RECT 100.095 80.150 100.355 80.410 ;
        RECT 100.415 80.150 100.675 80.410 ;
        RECT 121.330 80.150 121.590 80.410 ;
        RECT 121.650 80.150 121.910 80.410 ;
        RECT 121.970 80.150 122.230 80.410 ;
        RECT 122.290 80.150 122.550 80.410 ;
        RECT 122.610 80.150 122.870 80.410 ;
        RECT 143.525 80.150 143.785 80.410 ;
        RECT 143.845 80.150 144.105 80.410 ;
        RECT 144.165 80.150 144.425 80.410 ;
        RECT 144.485 80.150 144.745 80.410 ;
        RECT 144.805 80.150 145.065 80.410 ;
        RECT 76.940 74.710 77.200 74.970 ;
        RECT 77.260 74.710 77.520 74.970 ;
        RECT 77.580 74.710 77.840 74.970 ;
        RECT 77.900 74.710 78.160 74.970 ;
        RECT 78.220 74.710 78.480 74.970 ;
        RECT 99.135 74.710 99.395 74.970 ;
        RECT 99.455 74.710 99.715 74.970 ;
        RECT 99.775 74.710 100.035 74.970 ;
        RECT 100.095 74.710 100.355 74.970 ;
        RECT 100.415 74.710 100.675 74.970 ;
        RECT 121.330 74.710 121.590 74.970 ;
        RECT 121.650 74.710 121.910 74.970 ;
        RECT 121.970 74.710 122.230 74.970 ;
        RECT 122.290 74.710 122.550 74.970 ;
        RECT 122.610 74.710 122.870 74.970 ;
        RECT 143.525 74.710 143.785 74.970 ;
        RECT 143.845 74.710 144.105 74.970 ;
        RECT 144.165 74.710 144.425 74.970 ;
        RECT 144.485 74.710 144.745 74.970 ;
        RECT 144.805 74.710 145.065 74.970 ;
        RECT 76.940 69.270 77.200 69.530 ;
        RECT 77.260 69.270 77.520 69.530 ;
        RECT 77.580 69.270 77.840 69.530 ;
        RECT 77.900 69.270 78.160 69.530 ;
        RECT 78.220 69.270 78.480 69.530 ;
        RECT 99.135 69.270 99.395 69.530 ;
        RECT 99.455 69.270 99.715 69.530 ;
        RECT 99.775 69.270 100.035 69.530 ;
        RECT 100.095 69.270 100.355 69.530 ;
        RECT 100.415 69.270 100.675 69.530 ;
        RECT 121.330 69.270 121.590 69.530 ;
        RECT 121.650 69.270 121.910 69.530 ;
        RECT 121.970 69.270 122.230 69.530 ;
        RECT 122.290 69.270 122.550 69.530 ;
        RECT 122.610 69.270 122.870 69.530 ;
        RECT 143.525 69.270 143.785 69.530 ;
        RECT 143.845 69.270 144.105 69.530 ;
        RECT 144.165 69.270 144.425 69.530 ;
        RECT 144.485 69.270 144.745 69.530 ;
        RECT 144.805 69.270 145.065 69.530 ;
        RECT 76.940 63.830 77.200 64.090 ;
        RECT 77.260 63.830 77.520 64.090 ;
        RECT 77.580 63.830 77.840 64.090 ;
        RECT 77.900 63.830 78.160 64.090 ;
        RECT 78.220 63.830 78.480 64.090 ;
        RECT 99.135 63.830 99.395 64.090 ;
        RECT 99.455 63.830 99.715 64.090 ;
        RECT 99.775 63.830 100.035 64.090 ;
        RECT 100.095 63.830 100.355 64.090 ;
        RECT 100.415 63.830 100.675 64.090 ;
        RECT 121.330 63.830 121.590 64.090 ;
        RECT 121.650 63.830 121.910 64.090 ;
        RECT 121.970 63.830 122.230 64.090 ;
        RECT 122.290 63.830 122.550 64.090 ;
        RECT 122.610 63.830 122.870 64.090 ;
        RECT 143.525 63.830 143.785 64.090 ;
        RECT 143.845 63.830 144.105 64.090 ;
        RECT 144.165 63.830 144.425 64.090 ;
        RECT 144.485 63.830 144.745 64.090 ;
        RECT 144.805 63.830 145.065 64.090 ;
        RECT 76.940 58.390 77.200 58.650 ;
        RECT 77.260 58.390 77.520 58.650 ;
        RECT 77.580 58.390 77.840 58.650 ;
        RECT 77.900 58.390 78.160 58.650 ;
        RECT 78.220 58.390 78.480 58.650 ;
        RECT 99.135 58.390 99.395 58.650 ;
        RECT 99.455 58.390 99.715 58.650 ;
        RECT 99.775 58.390 100.035 58.650 ;
        RECT 100.095 58.390 100.355 58.650 ;
        RECT 100.415 58.390 100.675 58.650 ;
        RECT 121.330 58.390 121.590 58.650 ;
        RECT 121.650 58.390 121.910 58.650 ;
        RECT 121.970 58.390 122.230 58.650 ;
        RECT 122.290 58.390 122.550 58.650 ;
        RECT 122.610 58.390 122.870 58.650 ;
        RECT 143.525 58.390 143.785 58.650 ;
        RECT 143.845 58.390 144.105 58.650 ;
        RECT 144.165 58.390 144.425 58.650 ;
        RECT 144.485 58.390 144.745 58.650 ;
        RECT 144.805 58.390 145.065 58.650 ;
        RECT 76.940 52.950 77.200 53.210 ;
        RECT 77.260 52.950 77.520 53.210 ;
        RECT 77.580 52.950 77.840 53.210 ;
        RECT 77.900 52.950 78.160 53.210 ;
        RECT 78.220 52.950 78.480 53.210 ;
        RECT 99.135 52.950 99.395 53.210 ;
        RECT 99.455 52.950 99.715 53.210 ;
        RECT 99.775 52.950 100.035 53.210 ;
        RECT 100.095 52.950 100.355 53.210 ;
        RECT 100.415 52.950 100.675 53.210 ;
        RECT 121.330 52.950 121.590 53.210 ;
        RECT 121.650 52.950 121.910 53.210 ;
        RECT 121.970 52.950 122.230 53.210 ;
        RECT 122.290 52.950 122.550 53.210 ;
        RECT 122.610 52.950 122.870 53.210 ;
        RECT 143.525 52.950 143.785 53.210 ;
        RECT 143.845 52.950 144.105 53.210 ;
        RECT 144.165 52.950 144.425 53.210 ;
        RECT 144.485 52.950 144.745 53.210 ;
        RECT 144.805 52.950 145.065 53.210 ;
        RECT 76.940 47.510 77.200 47.770 ;
        RECT 77.260 47.510 77.520 47.770 ;
        RECT 77.580 47.510 77.840 47.770 ;
        RECT 77.900 47.510 78.160 47.770 ;
        RECT 78.220 47.510 78.480 47.770 ;
        RECT 99.135 47.510 99.395 47.770 ;
        RECT 99.455 47.510 99.715 47.770 ;
        RECT 99.775 47.510 100.035 47.770 ;
        RECT 100.095 47.510 100.355 47.770 ;
        RECT 100.415 47.510 100.675 47.770 ;
        RECT 121.330 47.510 121.590 47.770 ;
        RECT 121.650 47.510 121.910 47.770 ;
        RECT 121.970 47.510 122.230 47.770 ;
        RECT 122.290 47.510 122.550 47.770 ;
        RECT 122.610 47.510 122.870 47.770 ;
        RECT 143.525 47.510 143.785 47.770 ;
        RECT 143.845 47.510 144.105 47.770 ;
        RECT 144.165 47.510 144.425 47.770 ;
        RECT 144.485 47.510 144.745 47.770 ;
        RECT 144.805 47.510 145.065 47.770 ;
        RECT 76.940 42.070 77.200 42.330 ;
        RECT 77.260 42.070 77.520 42.330 ;
        RECT 77.580 42.070 77.840 42.330 ;
        RECT 77.900 42.070 78.160 42.330 ;
        RECT 78.220 42.070 78.480 42.330 ;
        RECT 99.135 42.070 99.395 42.330 ;
        RECT 99.455 42.070 99.715 42.330 ;
        RECT 99.775 42.070 100.035 42.330 ;
        RECT 100.095 42.070 100.355 42.330 ;
        RECT 100.415 42.070 100.675 42.330 ;
        RECT 121.330 42.070 121.590 42.330 ;
        RECT 121.650 42.070 121.910 42.330 ;
        RECT 121.970 42.070 122.230 42.330 ;
        RECT 122.290 42.070 122.550 42.330 ;
        RECT 122.610 42.070 122.870 42.330 ;
        RECT 143.525 42.070 143.785 42.330 ;
        RECT 143.845 42.070 144.105 42.330 ;
        RECT 144.165 42.070 144.425 42.330 ;
        RECT 144.485 42.070 144.745 42.330 ;
        RECT 144.805 42.070 145.065 42.330 ;
        RECT 76.940 36.630 77.200 36.890 ;
        RECT 77.260 36.630 77.520 36.890 ;
        RECT 77.580 36.630 77.840 36.890 ;
        RECT 77.900 36.630 78.160 36.890 ;
        RECT 78.220 36.630 78.480 36.890 ;
        RECT 99.135 36.630 99.395 36.890 ;
        RECT 99.455 36.630 99.715 36.890 ;
        RECT 99.775 36.630 100.035 36.890 ;
        RECT 100.095 36.630 100.355 36.890 ;
        RECT 100.415 36.630 100.675 36.890 ;
        RECT 121.330 36.630 121.590 36.890 ;
        RECT 121.650 36.630 121.910 36.890 ;
        RECT 121.970 36.630 122.230 36.890 ;
        RECT 122.290 36.630 122.550 36.890 ;
        RECT 122.610 36.630 122.870 36.890 ;
        RECT 143.525 36.630 143.785 36.890 ;
        RECT 143.845 36.630 144.105 36.890 ;
        RECT 144.165 36.630 144.425 36.890 ;
        RECT 144.485 36.630 144.745 36.890 ;
        RECT 144.805 36.630 145.065 36.890 ;
        RECT 76.940 31.190 77.200 31.450 ;
        RECT 77.260 31.190 77.520 31.450 ;
        RECT 77.580 31.190 77.840 31.450 ;
        RECT 77.900 31.190 78.160 31.450 ;
        RECT 78.220 31.190 78.480 31.450 ;
        RECT 99.135 31.190 99.395 31.450 ;
        RECT 99.455 31.190 99.715 31.450 ;
        RECT 99.775 31.190 100.035 31.450 ;
        RECT 100.095 31.190 100.355 31.450 ;
        RECT 100.415 31.190 100.675 31.450 ;
        RECT 121.330 31.190 121.590 31.450 ;
        RECT 121.650 31.190 121.910 31.450 ;
        RECT 121.970 31.190 122.230 31.450 ;
        RECT 122.290 31.190 122.550 31.450 ;
        RECT 122.610 31.190 122.870 31.450 ;
        RECT 143.525 31.190 143.785 31.450 ;
        RECT 143.845 31.190 144.105 31.450 ;
        RECT 144.165 31.190 144.425 31.450 ;
        RECT 144.485 31.190 144.745 31.450 ;
        RECT 144.805 31.190 145.065 31.450 ;
        RECT 76.940 25.750 77.200 26.010 ;
        RECT 77.260 25.750 77.520 26.010 ;
        RECT 77.580 25.750 77.840 26.010 ;
        RECT 77.900 25.750 78.160 26.010 ;
        RECT 78.220 25.750 78.480 26.010 ;
        RECT 99.135 25.750 99.395 26.010 ;
        RECT 99.455 25.750 99.715 26.010 ;
        RECT 99.775 25.750 100.035 26.010 ;
        RECT 100.095 25.750 100.355 26.010 ;
        RECT 100.415 25.750 100.675 26.010 ;
        RECT 121.330 25.750 121.590 26.010 ;
        RECT 121.650 25.750 121.910 26.010 ;
        RECT 121.970 25.750 122.230 26.010 ;
        RECT 122.290 25.750 122.550 26.010 ;
        RECT 122.610 25.750 122.870 26.010 ;
        RECT 143.525 25.750 143.785 26.010 ;
        RECT 143.845 25.750 144.105 26.010 ;
        RECT 144.165 25.750 144.425 26.010 ;
        RECT 144.485 25.750 144.745 26.010 ;
        RECT 144.805 25.750 145.065 26.010 ;
      LAYER met2 ;
        RECT 76.940 101.855 78.480 102.225 ;
        RECT 99.135 101.855 100.675 102.225 ;
        RECT 121.330 101.855 122.870 102.225 ;
        RECT 143.525 101.855 145.065 102.225 ;
        RECT 76.940 96.415 78.480 96.785 ;
        RECT 99.135 96.415 100.675 96.785 ;
        RECT 121.330 96.415 122.870 96.785 ;
        RECT 143.525 96.415 145.065 96.785 ;
        RECT 76.940 90.975 78.480 91.345 ;
        RECT 99.135 90.975 100.675 91.345 ;
        RECT 121.330 90.975 122.870 91.345 ;
        RECT 143.525 90.975 145.065 91.345 ;
        RECT 76.940 85.535 78.480 85.905 ;
        RECT 99.135 85.535 100.675 85.905 ;
        RECT 121.330 85.535 122.870 85.905 ;
        RECT 143.525 85.535 145.065 85.905 ;
        RECT 76.940 80.095 78.480 80.465 ;
        RECT 99.135 80.095 100.675 80.465 ;
        RECT 121.330 80.095 122.870 80.465 ;
        RECT 143.525 80.095 145.065 80.465 ;
        RECT 76.940 74.655 78.480 75.025 ;
        RECT 99.135 74.655 100.675 75.025 ;
        RECT 121.330 74.655 122.870 75.025 ;
        RECT 143.525 74.655 145.065 75.025 ;
        RECT 76.940 69.215 78.480 69.585 ;
        RECT 99.135 69.215 100.675 69.585 ;
        RECT 121.330 69.215 122.870 69.585 ;
        RECT 143.525 69.215 145.065 69.585 ;
        RECT 76.940 63.775 78.480 64.145 ;
        RECT 99.135 63.775 100.675 64.145 ;
        RECT 121.330 63.775 122.870 64.145 ;
        RECT 143.525 63.775 145.065 64.145 ;
        RECT 76.940 58.335 78.480 58.705 ;
        RECT 99.135 58.335 100.675 58.705 ;
        RECT 121.330 58.335 122.870 58.705 ;
        RECT 143.525 58.335 145.065 58.705 ;
        RECT 76.940 52.895 78.480 53.265 ;
        RECT 99.135 52.895 100.675 53.265 ;
        RECT 121.330 52.895 122.870 53.265 ;
        RECT 143.525 52.895 145.065 53.265 ;
        RECT 76.940 47.455 78.480 47.825 ;
        RECT 99.135 47.455 100.675 47.825 ;
        RECT 121.330 47.455 122.870 47.825 ;
        RECT 143.525 47.455 145.065 47.825 ;
        RECT 76.940 42.015 78.480 42.385 ;
        RECT 99.135 42.015 100.675 42.385 ;
        RECT 121.330 42.015 122.870 42.385 ;
        RECT 143.525 42.015 145.065 42.385 ;
        RECT 76.940 36.575 78.480 36.945 ;
        RECT 99.135 36.575 100.675 36.945 ;
        RECT 121.330 36.575 122.870 36.945 ;
        RECT 143.525 36.575 145.065 36.945 ;
        RECT 76.940 31.135 78.480 31.505 ;
        RECT 99.135 31.135 100.675 31.505 ;
        RECT 121.330 31.135 122.870 31.505 ;
        RECT 143.525 31.135 145.065 31.505 ;
        RECT 76.940 25.695 78.480 26.065 ;
        RECT 99.135 25.695 100.675 26.065 ;
        RECT 121.330 25.695 122.870 26.065 ;
        RECT 143.525 25.695 145.065 26.065 ;
      LAYER via2 ;
        RECT 76.970 101.900 77.250 102.180 ;
        RECT 77.370 101.900 77.650 102.180 ;
        RECT 77.770 101.900 78.050 102.180 ;
        RECT 78.170 101.900 78.450 102.180 ;
        RECT 99.165 101.900 99.445 102.180 ;
        RECT 99.565 101.900 99.845 102.180 ;
        RECT 99.965 101.900 100.245 102.180 ;
        RECT 100.365 101.900 100.645 102.180 ;
        RECT 121.360 101.900 121.640 102.180 ;
        RECT 121.760 101.900 122.040 102.180 ;
        RECT 122.160 101.900 122.440 102.180 ;
        RECT 122.560 101.900 122.840 102.180 ;
        RECT 143.555 101.900 143.835 102.180 ;
        RECT 143.955 101.900 144.235 102.180 ;
        RECT 144.355 101.900 144.635 102.180 ;
        RECT 144.755 101.900 145.035 102.180 ;
        RECT 76.970 96.460 77.250 96.740 ;
        RECT 77.370 96.460 77.650 96.740 ;
        RECT 77.770 96.460 78.050 96.740 ;
        RECT 78.170 96.460 78.450 96.740 ;
        RECT 99.165 96.460 99.445 96.740 ;
        RECT 99.565 96.460 99.845 96.740 ;
        RECT 99.965 96.460 100.245 96.740 ;
        RECT 100.365 96.460 100.645 96.740 ;
        RECT 121.360 96.460 121.640 96.740 ;
        RECT 121.760 96.460 122.040 96.740 ;
        RECT 122.160 96.460 122.440 96.740 ;
        RECT 122.560 96.460 122.840 96.740 ;
        RECT 143.555 96.460 143.835 96.740 ;
        RECT 143.955 96.460 144.235 96.740 ;
        RECT 144.355 96.460 144.635 96.740 ;
        RECT 144.755 96.460 145.035 96.740 ;
        RECT 76.970 91.020 77.250 91.300 ;
        RECT 77.370 91.020 77.650 91.300 ;
        RECT 77.770 91.020 78.050 91.300 ;
        RECT 78.170 91.020 78.450 91.300 ;
        RECT 99.165 91.020 99.445 91.300 ;
        RECT 99.565 91.020 99.845 91.300 ;
        RECT 99.965 91.020 100.245 91.300 ;
        RECT 100.365 91.020 100.645 91.300 ;
        RECT 121.360 91.020 121.640 91.300 ;
        RECT 121.760 91.020 122.040 91.300 ;
        RECT 122.160 91.020 122.440 91.300 ;
        RECT 122.560 91.020 122.840 91.300 ;
        RECT 143.555 91.020 143.835 91.300 ;
        RECT 143.955 91.020 144.235 91.300 ;
        RECT 144.355 91.020 144.635 91.300 ;
        RECT 144.755 91.020 145.035 91.300 ;
        RECT 76.970 85.580 77.250 85.860 ;
        RECT 77.370 85.580 77.650 85.860 ;
        RECT 77.770 85.580 78.050 85.860 ;
        RECT 78.170 85.580 78.450 85.860 ;
        RECT 99.165 85.580 99.445 85.860 ;
        RECT 99.565 85.580 99.845 85.860 ;
        RECT 99.965 85.580 100.245 85.860 ;
        RECT 100.365 85.580 100.645 85.860 ;
        RECT 121.360 85.580 121.640 85.860 ;
        RECT 121.760 85.580 122.040 85.860 ;
        RECT 122.160 85.580 122.440 85.860 ;
        RECT 122.560 85.580 122.840 85.860 ;
        RECT 143.555 85.580 143.835 85.860 ;
        RECT 143.955 85.580 144.235 85.860 ;
        RECT 144.355 85.580 144.635 85.860 ;
        RECT 144.755 85.580 145.035 85.860 ;
        RECT 76.970 80.140 77.250 80.420 ;
        RECT 77.370 80.140 77.650 80.420 ;
        RECT 77.770 80.140 78.050 80.420 ;
        RECT 78.170 80.140 78.450 80.420 ;
        RECT 99.165 80.140 99.445 80.420 ;
        RECT 99.565 80.140 99.845 80.420 ;
        RECT 99.965 80.140 100.245 80.420 ;
        RECT 100.365 80.140 100.645 80.420 ;
        RECT 121.360 80.140 121.640 80.420 ;
        RECT 121.760 80.140 122.040 80.420 ;
        RECT 122.160 80.140 122.440 80.420 ;
        RECT 122.560 80.140 122.840 80.420 ;
        RECT 143.555 80.140 143.835 80.420 ;
        RECT 143.955 80.140 144.235 80.420 ;
        RECT 144.355 80.140 144.635 80.420 ;
        RECT 144.755 80.140 145.035 80.420 ;
        RECT 76.970 74.700 77.250 74.980 ;
        RECT 77.370 74.700 77.650 74.980 ;
        RECT 77.770 74.700 78.050 74.980 ;
        RECT 78.170 74.700 78.450 74.980 ;
        RECT 99.165 74.700 99.445 74.980 ;
        RECT 99.565 74.700 99.845 74.980 ;
        RECT 99.965 74.700 100.245 74.980 ;
        RECT 100.365 74.700 100.645 74.980 ;
        RECT 121.360 74.700 121.640 74.980 ;
        RECT 121.760 74.700 122.040 74.980 ;
        RECT 122.160 74.700 122.440 74.980 ;
        RECT 122.560 74.700 122.840 74.980 ;
        RECT 143.555 74.700 143.835 74.980 ;
        RECT 143.955 74.700 144.235 74.980 ;
        RECT 144.355 74.700 144.635 74.980 ;
        RECT 144.755 74.700 145.035 74.980 ;
        RECT 76.970 69.260 77.250 69.540 ;
        RECT 77.370 69.260 77.650 69.540 ;
        RECT 77.770 69.260 78.050 69.540 ;
        RECT 78.170 69.260 78.450 69.540 ;
        RECT 99.165 69.260 99.445 69.540 ;
        RECT 99.565 69.260 99.845 69.540 ;
        RECT 99.965 69.260 100.245 69.540 ;
        RECT 100.365 69.260 100.645 69.540 ;
        RECT 121.360 69.260 121.640 69.540 ;
        RECT 121.760 69.260 122.040 69.540 ;
        RECT 122.160 69.260 122.440 69.540 ;
        RECT 122.560 69.260 122.840 69.540 ;
        RECT 143.555 69.260 143.835 69.540 ;
        RECT 143.955 69.260 144.235 69.540 ;
        RECT 144.355 69.260 144.635 69.540 ;
        RECT 144.755 69.260 145.035 69.540 ;
        RECT 76.970 63.820 77.250 64.100 ;
        RECT 77.370 63.820 77.650 64.100 ;
        RECT 77.770 63.820 78.050 64.100 ;
        RECT 78.170 63.820 78.450 64.100 ;
        RECT 99.165 63.820 99.445 64.100 ;
        RECT 99.565 63.820 99.845 64.100 ;
        RECT 99.965 63.820 100.245 64.100 ;
        RECT 100.365 63.820 100.645 64.100 ;
        RECT 121.360 63.820 121.640 64.100 ;
        RECT 121.760 63.820 122.040 64.100 ;
        RECT 122.160 63.820 122.440 64.100 ;
        RECT 122.560 63.820 122.840 64.100 ;
        RECT 143.555 63.820 143.835 64.100 ;
        RECT 143.955 63.820 144.235 64.100 ;
        RECT 144.355 63.820 144.635 64.100 ;
        RECT 144.755 63.820 145.035 64.100 ;
        RECT 76.970 58.380 77.250 58.660 ;
        RECT 77.370 58.380 77.650 58.660 ;
        RECT 77.770 58.380 78.050 58.660 ;
        RECT 78.170 58.380 78.450 58.660 ;
        RECT 99.165 58.380 99.445 58.660 ;
        RECT 99.565 58.380 99.845 58.660 ;
        RECT 99.965 58.380 100.245 58.660 ;
        RECT 100.365 58.380 100.645 58.660 ;
        RECT 121.360 58.380 121.640 58.660 ;
        RECT 121.760 58.380 122.040 58.660 ;
        RECT 122.160 58.380 122.440 58.660 ;
        RECT 122.560 58.380 122.840 58.660 ;
        RECT 143.555 58.380 143.835 58.660 ;
        RECT 143.955 58.380 144.235 58.660 ;
        RECT 144.355 58.380 144.635 58.660 ;
        RECT 144.755 58.380 145.035 58.660 ;
        RECT 76.970 52.940 77.250 53.220 ;
        RECT 77.370 52.940 77.650 53.220 ;
        RECT 77.770 52.940 78.050 53.220 ;
        RECT 78.170 52.940 78.450 53.220 ;
        RECT 99.165 52.940 99.445 53.220 ;
        RECT 99.565 52.940 99.845 53.220 ;
        RECT 99.965 52.940 100.245 53.220 ;
        RECT 100.365 52.940 100.645 53.220 ;
        RECT 121.360 52.940 121.640 53.220 ;
        RECT 121.760 52.940 122.040 53.220 ;
        RECT 122.160 52.940 122.440 53.220 ;
        RECT 122.560 52.940 122.840 53.220 ;
        RECT 143.555 52.940 143.835 53.220 ;
        RECT 143.955 52.940 144.235 53.220 ;
        RECT 144.355 52.940 144.635 53.220 ;
        RECT 144.755 52.940 145.035 53.220 ;
        RECT 76.970 47.500 77.250 47.780 ;
        RECT 77.370 47.500 77.650 47.780 ;
        RECT 77.770 47.500 78.050 47.780 ;
        RECT 78.170 47.500 78.450 47.780 ;
        RECT 99.165 47.500 99.445 47.780 ;
        RECT 99.565 47.500 99.845 47.780 ;
        RECT 99.965 47.500 100.245 47.780 ;
        RECT 100.365 47.500 100.645 47.780 ;
        RECT 121.360 47.500 121.640 47.780 ;
        RECT 121.760 47.500 122.040 47.780 ;
        RECT 122.160 47.500 122.440 47.780 ;
        RECT 122.560 47.500 122.840 47.780 ;
        RECT 143.555 47.500 143.835 47.780 ;
        RECT 143.955 47.500 144.235 47.780 ;
        RECT 144.355 47.500 144.635 47.780 ;
        RECT 144.755 47.500 145.035 47.780 ;
        RECT 76.970 42.060 77.250 42.340 ;
        RECT 77.370 42.060 77.650 42.340 ;
        RECT 77.770 42.060 78.050 42.340 ;
        RECT 78.170 42.060 78.450 42.340 ;
        RECT 99.165 42.060 99.445 42.340 ;
        RECT 99.565 42.060 99.845 42.340 ;
        RECT 99.965 42.060 100.245 42.340 ;
        RECT 100.365 42.060 100.645 42.340 ;
        RECT 121.360 42.060 121.640 42.340 ;
        RECT 121.760 42.060 122.040 42.340 ;
        RECT 122.160 42.060 122.440 42.340 ;
        RECT 122.560 42.060 122.840 42.340 ;
        RECT 143.555 42.060 143.835 42.340 ;
        RECT 143.955 42.060 144.235 42.340 ;
        RECT 144.355 42.060 144.635 42.340 ;
        RECT 144.755 42.060 145.035 42.340 ;
        RECT 76.970 36.620 77.250 36.900 ;
        RECT 77.370 36.620 77.650 36.900 ;
        RECT 77.770 36.620 78.050 36.900 ;
        RECT 78.170 36.620 78.450 36.900 ;
        RECT 99.165 36.620 99.445 36.900 ;
        RECT 99.565 36.620 99.845 36.900 ;
        RECT 99.965 36.620 100.245 36.900 ;
        RECT 100.365 36.620 100.645 36.900 ;
        RECT 121.360 36.620 121.640 36.900 ;
        RECT 121.760 36.620 122.040 36.900 ;
        RECT 122.160 36.620 122.440 36.900 ;
        RECT 122.560 36.620 122.840 36.900 ;
        RECT 143.555 36.620 143.835 36.900 ;
        RECT 143.955 36.620 144.235 36.900 ;
        RECT 144.355 36.620 144.635 36.900 ;
        RECT 144.755 36.620 145.035 36.900 ;
        RECT 76.970 31.180 77.250 31.460 ;
        RECT 77.370 31.180 77.650 31.460 ;
        RECT 77.770 31.180 78.050 31.460 ;
        RECT 78.170 31.180 78.450 31.460 ;
        RECT 99.165 31.180 99.445 31.460 ;
        RECT 99.565 31.180 99.845 31.460 ;
        RECT 99.965 31.180 100.245 31.460 ;
        RECT 100.365 31.180 100.645 31.460 ;
        RECT 121.360 31.180 121.640 31.460 ;
        RECT 121.760 31.180 122.040 31.460 ;
        RECT 122.160 31.180 122.440 31.460 ;
        RECT 122.560 31.180 122.840 31.460 ;
        RECT 143.555 31.180 143.835 31.460 ;
        RECT 143.955 31.180 144.235 31.460 ;
        RECT 144.355 31.180 144.635 31.460 ;
        RECT 144.755 31.180 145.035 31.460 ;
        RECT 76.970 25.740 77.250 26.020 ;
        RECT 77.370 25.740 77.650 26.020 ;
        RECT 77.770 25.740 78.050 26.020 ;
        RECT 78.170 25.740 78.450 26.020 ;
        RECT 99.165 25.740 99.445 26.020 ;
        RECT 99.565 25.740 99.845 26.020 ;
        RECT 99.965 25.740 100.245 26.020 ;
        RECT 100.365 25.740 100.645 26.020 ;
        RECT 121.360 25.740 121.640 26.020 ;
        RECT 121.760 25.740 122.040 26.020 ;
        RECT 122.160 25.740 122.440 26.020 ;
        RECT 122.560 25.740 122.840 26.020 ;
        RECT 143.555 25.740 143.835 26.020 ;
        RECT 143.955 25.740 144.235 26.020 ;
        RECT 144.355 25.740 144.635 26.020 ;
        RECT 144.755 25.740 145.035 26.020 ;
      LAYER met3 ;
        RECT 76.920 101.875 78.500 102.205 ;
        RECT 99.115 101.875 100.695 102.205 ;
        RECT 121.310 101.875 122.890 102.205 ;
        RECT 143.505 101.875 145.085 102.205 ;
        RECT 76.920 96.435 78.500 96.765 ;
        RECT 99.115 96.435 100.695 96.765 ;
        RECT 121.310 96.435 122.890 96.765 ;
        RECT 143.505 96.435 145.085 96.765 ;
        RECT 76.920 90.995 78.500 91.325 ;
        RECT 99.115 90.995 100.695 91.325 ;
        RECT 121.310 90.995 122.890 91.325 ;
        RECT 143.505 90.995 145.085 91.325 ;
        RECT 76.920 85.555 78.500 85.885 ;
        RECT 99.115 85.555 100.695 85.885 ;
        RECT 121.310 85.555 122.890 85.885 ;
        RECT 143.505 85.555 145.085 85.885 ;
        RECT 76.920 80.115 78.500 80.445 ;
        RECT 99.115 80.115 100.695 80.445 ;
        RECT 121.310 80.115 122.890 80.445 ;
        RECT 143.505 80.115 145.085 80.445 ;
        RECT 76.920 74.675 78.500 75.005 ;
        RECT 99.115 74.675 100.695 75.005 ;
        RECT 121.310 74.675 122.890 75.005 ;
        RECT 143.505 74.675 145.085 75.005 ;
        RECT 76.920 69.235 78.500 69.565 ;
        RECT 99.115 69.235 100.695 69.565 ;
        RECT 121.310 69.235 122.890 69.565 ;
        RECT 143.505 69.235 145.085 69.565 ;
        RECT 76.920 63.795 78.500 64.125 ;
        RECT 99.115 63.795 100.695 64.125 ;
        RECT 121.310 63.795 122.890 64.125 ;
        RECT 143.505 63.795 145.085 64.125 ;
        RECT 76.920 58.355 78.500 58.685 ;
        RECT 99.115 58.355 100.695 58.685 ;
        RECT 121.310 58.355 122.890 58.685 ;
        RECT 143.505 58.355 145.085 58.685 ;
        RECT 76.920 52.915 78.500 53.245 ;
        RECT 99.115 52.915 100.695 53.245 ;
        RECT 121.310 52.915 122.890 53.245 ;
        RECT 143.505 52.915 145.085 53.245 ;
        RECT 76.920 47.475 78.500 47.805 ;
        RECT 99.115 47.475 100.695 47.805 ;
        RECT 121.310 47.475 122.890 47.805 ;
        RECT 143.505 47.475 145.085 47.805 ;
        RECT 76.920 42.035 78.500 42.365 ;
        RECT 99.115 42.035 100.695 42.365 ;
        RECT 121.310 42.035 122.890 42.365 ;
        RECT 143.505 42.035 145.085 42.365 ;
        RECT 76.920 36.595 78.500 36.925 ;
        RECT 99.115 36.595 100.695 36.925 ;
        RECT 121.310 36.595 122.890 36.925 ;
        RECT 143.505 36.595 145.085 36.925 ;
        RECT 76.920 31.155 78.500 31.485 ;
        RECT 99.115 31.155 100.695 31.485 ;
        RECT 121.310 31.155 122.890 31.485 ;
        RECT 143.505 31.155 145.085 31.485 ;
        RECT 76.920 25.715 78.500 26.045 ;
        RECT 99.115 25.715 100.695 26.045 ;
        RECT 121.310 25.715 122.890 26.045 ;
        RECT 143.505 25.715 145.085 26.045 ;
      LAYER via3 ;
        RECT 76.950 101.880 77.270 102.200 ;
        RECT 77.350 101.880 77.670 102.200 ;
        RECT 77.750 101.880 78.070 102.200 ;
        RECT 78.150 101.880 78.470 102.200 ;
        RECT 99.145 101.880 99.465 102.200 ;
        RECT 99.545 101.880 99.865 102.200 ;
        RECT 99.945 101.880 100.265 102.200 ;
        RECT 100.345 101.880 100.665 102.200 ;
        RECT 121.340 101.880 121.660 102.200 ;
        RECT 121.740 101.880 122.060 102.200 ;
        RECT 122.140 101.880 122.460 102.200 ;
        RECT 122.540 101.880 122.860 102.200 ;
        RECT 143.535 101.880 143.855 102.200 ;
        RECT 143.935 101.880 144.255 102.200 ;
        RECT 144.335 101.880 144.655 102.200 ;
        RECT 144.735 101.880 145.055 102.200 ;
        RECT 76.950 96.440 77.270 96.760 ;
        RECT 77.350 96.440 77.670 96.760 ;
        RECT 77.750 96.440 78.070 96.760 ;
        RECT 78.150 96.440 78.470 96.760 ;
        RECT 99.145 96.440 99.465 96.760 ;
        RECT 99.545 96.440 99.865 96.760 ;
        RECT 99.945 96.440 100.265 96.760 ;
        RECT 100.345 96.440 100.665 96.760 ;
        RECT 121.340 96.440 121.660 96.760 ;
        RECT 121.740 96.440 122.060 96.760 ;
        RECT 122.140 96.440 122.460 96.760 ;
        RECT 122.540 96.440 122.860 96.760 ;
        RECT 143.535 96.440 143.855 96.760 ;
        RECT 143.935 96.440 144.255 96.760 ;
        RECT 144.335 96.440 144.655 96.760 ;
        RECT 144.735 96.440 145.055 96.760 ;
        RECT 76.950 91.000 77.270 91.320 ;
        RECT 77.350 91.000 77.670 91.320 ;
        RECT 77.750 91.000 78.070 91.320 ;
        RECT 78.150 91.000 78.470 91.320 ;
        RECT 99.145 91.000 99.465 91.320 ;
        RECT 99.545 91.000 99.865 91.320 ;
        RECT 99.945 91.000 100.265 91.320 ;
        RECT 100.345 91.000 100.665 91.320 ;
        RECT 121.340 91.000 121.660 91.320 ;
        RECT 121.740 91.000 122.060 91.320 ;
        RECT 122.140 91.000 122.460 91.320 ;
        RECT 122.540 91.000 122.860 91.320 ;
        RECT 143.535 91.000 143.855 91.320 ;
        RECT 143.935 91.000 144.255 91.320 ;
        RECT 144.335 91.000 144.655 91.320 ;
        RECT 144.735 91.000 145.055 91.320 ;
        RECT 76.950 85.560 77.270 85.880 ;
        RECT 77.350 85.560 77.670 85.880 ;
        RECT 77.750 85.560 78.070 85.880 ;
        RECT 78.150 85.560 78.470 85.880 ;
        RECT 99.145 85.560 99.465 85.880 ;
        RECT 99.545 85.560 99.865 85.880 ;
        RECT 99.945 85.560 100.265 85.880 ;
        RECT 100.345 85.560 100.665 85.880 ;
        RECT 121.340 85.560 121.660 85.880 ;
        RECT 121.740 85.560 122.060 85.880 ;
        RECT 122.140 85.560 122.460 85.880 ;
        RECT 122.540 85.560 122.860 85.880 ;
        RECT 143.535 85.560 143.855 85.880 ;
        RECT 143.935 85.560 144.255 85.880 ;
        RECT 144.335 85.560 144.655 85.880 ;
        RECT 144.735 85.560 145.055 85.880 ;
        RECT 76.950 80.120 77.270 80.440 ;
        RECT 77.350 80.120 77.670 80.440 ;
        RECT 77.750 80.120 78.070 80.440 ;
        RECT 78.150 80.120 78.470 80.440 ;
        RECT 99.145 80.120 99.465 80.440 ;
        RECT 99.545 80.120 99.865 80.440 ;
        RECT 99.945 80.120 100.265 80.440 ;
        RECT 100.345 80.120 100.665 80.440 ;
        RECT 121.340 80.120 121.660 80.440 ;
        RECT 121.740 80.120 122.060 80.440 ;
        RECT 122.140 80.120 122.460 80.440 ;
        RECT 122.540 80.120 122.860 80.440 ;
        RECT 143.535 80.120 143.855 80.440 ;
        RECT 143.935 80.120 144.255 80.440 ;
        RECT 144.335 80.120 144.655 80.440 ;
        RECT 144.735 80.120 145.055 80.440 ;
        RECT 76.950 74.680 77.270 75.000 ;
        RECT 77.350 74.680 77.670 75.000 ;
        RECT 77.750 74.680 78.070 75.000 ;
        RECT 78.150 74.680 78.470 75.000 ;
        RECT 99.145 74.680 99.465 75.000 ;
        RECT 99.545 74.680 99.865 75.000 ;
        RECT 99.945 74.680 100.265 75.000 ;
        RECT 100.345 74.680 100.665 75.000 ;
        RECT 121.340 74.680 121.660 75.000 ;
        RECT 121.740 74.680 122.060 75.000 ;
        RECT 122.140 74.680 122.460 75.000 ;
        RECT 122.540 74.680 122.860 75.000 ;
        RECT 143.535 74.680 143.855 75.000 ;
        RECT 143.935 74.680 144.255 75.000 ;
        RECT 144.335 74.680 144.655 75.000 ;
        RECT 144.735 74.680 145.055 75.000 ;
        RECT 76.950 69.240 77.270 69.560 ;
        RECT 77.350 69.240 77.670 69.560 ;
        RECT 77.750 69.240 78.070 69.560 ;
        RECT 78.150 69.240 78.470 69.560 ;
        RECT 99.145 69.240 99.465 69.560 ;
        RECT 99.545 69.240 99.865 69.560 ;
        RECT 99.945 69.240 100.265 69.560 ;
        RECT 100.345 69.240 100.665 69.560 ;
        RECT 121.340 69.240 121.660 69.560 ;
        RECT 121.740 69.240 122.060 69.560 ;
        RECT 122.140 69.240 122.460 69.560 ;
        RECT 122.540 69.240 122.860 69.560 ;
        RECT 143.535 69.240 143.855 69.560 ;
        RECT 143.935 69.240 144.255 69.560 ;
        RECT 144.335 69.240 144.655 69.560 ;
        RECT 144.735 69.240 145.055 69.560 ;
        RECT 76.950 63.800 77.270 64.120 ;
        RECT 77.350 63.800 77.670 64.120 ;
        RECT 77.750 63.800 78.070 64.120 ;
        RECT 78.150 63.800 78.470 64.120 ;
        RECT 99.145 63.800 99.465 64.120 ;
        RECT 99.545 63.800 99.865 64.120 ;
        RECT 99.945 63.800 100.265 64.120 ;
        RECT 100.345 63.800 100.665 64.120 ;
        RECT 121.340 63.800 121.660 64.120 ;
        RECT 121.740 63.800 122.060 64.120 ;
        RECT 122.140 63.800 122.460 64.120 ;
        RECT 122.540 63.800 122.860 64.120 ;
        RECT 143.535 63.800 143.855 64.120 ;
        RECT 143.935 63.800 144.255 64.120 ;
        RECT 144.335 63.800 144.655 64.120 ;
        RECT 144.735 63.800 145.055 64.120 ;
        RECT 76.950 58.360 77.270 58.680 ;
        RECT 77.350 58.360 77.670 58.680 ;
        RECT 77.750 58.360 78.070 58.680 ;
        RECT 78.150 58.360 78.470 58.680 ;
        RECT 99.145 58.360 99.465 58.680 ;
        RECT 99.545 58.360 99.865 58.680 ;
        RECT 99.945 58.360 100.265 58.680 ;
        RECT 100.345 58.360 100.665 58.680 ;
        RECT 121.340 58.360 121.660 58.680 ;
        RECT 121.740 58.360 122.060 58.680 ;
        RECT 122.140 58.360 122.460 58.680 ;
        RECT 122.540 58.360 122.860 58.680 ;
        RECT 143.535 58.360 143.855 58.680 ;
        RECT 143.935 58.360 144.255 58.680 ;
        RECT 144.335 58.360 144.655 58.680 ;
        RECT 144.735 58.360 145.055 58.680 ;
        RECT 76.950 52.920 77.270 53.240 ;
        RECT 77.350 52.920 77.670 53.240 ;
        RECT 77.750 52.920 78.070 53.240 ;
        RECT 78.150 52.920 78.470 53.240 ;
        RECT 99.145 52.920 99.465 53.240 ;
        RECT 99.545 52.920 99.865 53.240 ;
        RECT 99.945 52.920 100.265 53.240 ;
        RECT 100.345 52.920 100.665 53.240 ;
        RECT 121.340 52.920 121.660 53.240 ;
        RECT 121.740 52.920 122.060 53.240 ;
        RECT 122.140 52.920 122.460 53.240 ;
        RECT 122.540 52.920 122.860 53.240 ;
        RECT 143.535 52.920 143.855 53.240 ;
        RECT 143.935 52.920 144.255 53.240 ;
        RECT 144.335 52.920 144.655 53.240 ;
        RECT 144.735 52.920 145.055 53.240 ;
        RECT 76.950 47.480 77.270 47.800 ;
        RECT 77.350 47.480 77.670 47.800 ;
        RECT 77.750 47.480 78.070 47.800 ;
        RECT 78.150 47.480 78.470 47.800 ;
        RECT 99.145 47.480 99.465 47.800 ;
        RECT 99.545 47.480 99.865 47.800 ;
        RECT 99.945 47.480 100.265 47.800 ;
        RECT 100.345 47.480 100.665 47.800 ;
        RECT 121.340 47.480 121.660 47.800 ;
        RECT 121.740 47.480 122.060 47.800 ;
        RECT 122.140 47.480 122.460 47.800 ;
        RECT 122.540 47.480 122.860 47.800 ;
        RECT 143.535 47.480 143.855 47.800 ;
        RECT 143.935 47.480 144.255 47.800 ;
        RECT 144.335 47.480 144.655 47.800 ;
        RECT 144.735 47.480 145.055 47.800 ;
        RECT 76.950 42.040 77.270 42.360 ;
        RECT 77.350 42.040 77.670 42.360 ;
        RECT 77.750 42.040 78.070 42.360 ;
        RECT 78.150 42.040 78.470 42.360 ;
        RECT 99.145 42.040 99.465 42.360 ;
        RECT 99.545 42.040 99.865 42.360 ;
        RECT 99.945 42.040 100.265 42.360 ;
        RECT 100.345 42.040 100.665 42.360 ;
        RECT 121.340 42.040 121.660 42.360 ;
        RECT 121.740 42.040 122.060 42.360 ;
        RECT 122.140 42.040 122.460 42.360 ;
        RECT 122.540 42.040 122.860 42.360 ;
        RECT 143.535 42.040 143.855 42.360 ;
        RECT 143.935 42.040 144.255 42.360 ;
        RECT 144.335 42.040 144.655 42.360 ;
        RECT 144.735 42.040 145.055 42.360 ;
        RECT 76.950 36.600 77.270 36.920 ;
        RECT 77.350 36.600 77.670 36.920 ;
        RECT 77.750 36.600 78.070 36.920 ;
        RECT 78.150 36.600 78.470 36.920 ;
        RECT 99.145 36.600 99.465 36.920 ;
        RECT 99.545 36.600 99.865 36.920 ;
        RECT 99.945 36.600 100.265 36.920 ;
        RECT 100.345 36.600 100.665 36.920 ;
        RECT 121.340 36.600 121.660 36.920 ;
        RECT 121.740 36.600 122.060 36.920 ;
        RECT 122.140 36.600 122.460 36.920 ;
        RECT 122.540 36.600 122.860 36.920 ;
        RECT 143.535 36.600 143.855 36.920 ;
        RECT 143.935 36.600 144.255 36.920 ;
        RECT 144.335 36.600 144.655 36.920 ;
        RECT 144.735 36.600 145.055 36.920 ;
        RECT 76.950 31.160 77.270 31.480 ;
        RECT 77.350 31.160 77.670 31.480 ;
        RECT 77.750 31.160 78.070 31.480 ;
        RECT 78.150 31.160 78.470 31.480 ;
        RECT 99.145 31.160 99.465 31.480 ;
        RECT 99.545 31.160 99.865 31.480 ;
        RECT 99.945 31.160 100.265 31.480 ;
        RECT 100.345 31.160 100.665 31.480 ;
        RECT 121.340 31.160 121.660 31.480 ;
        RECT 121.740 31.160 122.060 31.480 ;
        RECT 122.140 31.160 122.460 31.480 ;
        RECT 122.540 31.160 122.860 31.480 ;
        RECT 143.535 31.160 143.855 31.480 ;
        RECT 143.935 31.160 144.255 31.480 ;
        RECT 144.335 31.160 144.655 31.480 ;
        RECT 144.735 31.160 145.055 31.480 ;
        RECT 76.950 25.720 77.270 26.040 ;
        RECT 77.350 25.720 77.670 26.040 ;
        RECT 77.750 25.720 78.070 26.040 ;
        RECT 78.150 25.720 78.470 26.040 ;
        RECT 99.145 25.720 99.465 26.040 ;
        RECT 99.545 25.720 99.865 26.040 ;
        RECT 99.945 25.720 100.265 26.040 ;
        RECT 100.345 25.720 100.665 26.040 ;
        RECT 121.340 25.720 121.660 26.040 ;
        RECT 121.740 25.720 122.060 26.040 ;
        RECT 122.140 25.720 122.460 26.040 ;
        RECT 122.540 25.720 122.860 26.040 ;
        RECT 143.535 25.720 143.855 26.040 ;
        RECT 143.935 25.720 144.255 26.040 ;
        RECT 144.335 25.720 144.655 26.040 ;
        RECT 144.735 25.720 145.055 26.040 ;
      LAYER met4 ;
        RECT 76.910 25.640 78.510 102.280 ;
        RECT 99.105 25.640 100.705 102.280 ;
        RECT 121.300 25.640 122.900 102.280 ;
        RECT 143.495 25.640 145.095 102.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN sky130_ef_sc_hd__decap_12_364/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 25.795 57.215 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_364/VNB
  PIN sky130_fd_sc_hd__decap_3_65/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 25.795 55.835 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_65/VNB
  PIN sky130_ef_sc_hd__decap_12_363/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 31.235 57.215 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_363/VNB
  PIN sky130_fd_sc_hd__decap_3_64/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 31.235 55.835 31.405 ;
    END
  END sky130_fd_sc_hd__decap_3_64/VNB
  PIN sky130_ef_sc_hd__decap_12_362/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 25.795 62.735 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_362/VNB
  PIN sky130_ef_sc_hd__decap_12_361/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 31.235 62.735 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_361/VNB
  PIN sky130_fd_sc_hd__fill_1_108/VNB
    PORT
      LAYER pwell ;
        RECT 68.080 25.825 68.200 25.935 ;
    END
  END sky130_fd_sc_hd__fill_1_108/VNB
  PIN sky130_ef_sc_hd__decap_12_360/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 25.795 69.175 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_360/VNB
  PIN sky130_ef_sc_hd__decap_12_359/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 31.375 68.255 31.405 ;
        RECT 68.080 31.265 68.255 31.375 ;
        RECT 68.085 31.235 68.255 31.265 ;
    END
  END sky130_ef_sc_hd__decap_12_359/VNB
  PIN sky130_ef_sc_hd__decap_12_358/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 25.795 74.695 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_358/VNB
  PIN sky130_ef_sc_hd__decap_12_357/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 31.235 73.775 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_357/VNB
  PIN sky130_fd_sc_hd__decap_4_10/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 31.235 79.295 31.405 ;
    END
  END sky130_fd_sc_hd__decap_4_10/VNB
  PIN sky130_fd_sc_hd__decap_3_63/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 25.795 80.215 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_63/VNB
  PIN sky130_ef_sc_hd__decap_12_356/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 25.795 82.055 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_356/VNB
  PIN sky130_fd_sc_hd__fill_1_107/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 31.265 81.080 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_107/VNB
  PIN sky130_ef_sc_hd__decap_12_355/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 31.235 82.055 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_355/VNB
  PIN sky130_ef_sc_hd__decap_12_354/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 25.795 87.575 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_354/VNB
  PIN sky130_ef_sc_hd__decap_12_353/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 31.235 87.575 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_353/VNB
  PIN sky130_fd_sc_hd__decap_3_62/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 25.795 93.095 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_62/VNB
  PIN sky130_ef_sc_hd__decap_12_352/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 25.795 94.935 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_352/VNB
  PIN sky130_ef_sc_hd__decap_12_351/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 31.235 93.095 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_351/VNB
  PIN sky130_ef_sc_hd__decap_12_350/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 25.795 100.455 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_350/VNB
  PIN sky130_ef_sc_hd__decap_12_349/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 31.235 98.615 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_349/VNB
  PIN sky130_fd_sc_hd__decap_3_61/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 25.795 105.975 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_61/VNB
  PIN sky130_ef_sc_hd__decap_12_348/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 25.795 107.815 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_348/VNB
  PIN sky130_fd_sc_hd__decap_6_55/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 31.235 104.135 31.405 ;
    END
  END sky130_fd_sc_hd__decap_6_55/VNB
  PIN sky130_fd_sc_hd__fill_1_106/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 31.265 106.840 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_106/VNB
  PIN sky130_ef_sc_hd__decap_12_347/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 31.235 107.815 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_347/VNB
  PIN sky130_ef_sc_hd__decap_12_346/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 25.795 113.335 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_346/VNB
  PIN sky130_ef_sc_hd__decap_12_345/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 31.235 113.335 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_345/VNB
  PIN sky130_fd_sc_hd__decap_3_60/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 25.795 118.855 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_60/VNB
  PIN sky130_ef_sc_hd__decap_12_343/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 31.235 118.855 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_343/VNB
  PIN sky130_ef_sc_hd__decap_12_344/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 25.795 120.695 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_344/VNB
  PIN sky130_ef_sc_hd__decap_12_342/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 25.795 126.215 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_342/VNB
  PIN sky130_ef_sc_hd__decap_12_341/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 31.235 124.375 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_341/VNB
  PIN sky130_fd_sc_hd__decap_3_59/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 25.795 131.735 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_59/VNB
  PIN sky130_fd_sc_hd__decap_6_54/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 31.235 129.895 31.405 ;
    END
  END sky130_fd_sc_hd__decap_6_54/VNB
  PIN sky130_fd_sc_hd__fill_1_105/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 31.265 132.600 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_105/VNB
  PIN sky130_ef_sc_hd__decap_12_340/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 25.795 133.575 25.965 ;
    END
  END sky130_ef_sc_hd__decap_12_340/VNB
  PIN sky130_ef_sc_hd__decap_12_339/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 31.235 133.575 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_339/VNB
  PIN sky130_fd_sc_hd__decap_8_19/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 25.795 139.095 25.965 ;
    END
  END sky130_fd_sc_hd__decap_8_19/VNB
  PIN sky130_fd_sc_hd__fill_1_104/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 25.825 142.720 25.935 ;
    END
  END sky130_fd_sc_hd__fill_1_104/VNB
  PIN sky130_fd_sc_hd__decap_8_18/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 31.235 139.095 31.405 ;
    END
  END sky130_fd_sc_hd__decap_8_18/VNB
  PIN sky130_fd_sc_hd__fill_1_103/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 31.265 142.720 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_103/VNB
  PIN sky130_fd_sc_hd__decap_3_58/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 25.795 144.155 25.965 ;
    END
  END sky130_fd_sc_hd__decap_3_58/VNB
  PIN sky130_fd_sc_hd__decap_3_57/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 31.235 144.155 31.405 ;
    END
  END sky130_fd_sc_hd__decap_3_57/VNB
  PIN sky130_ef_sc_hd__decap_12_336/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 31.235 69.175 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_336/VNB
  PIN sky130_ef_sc_hd__decap_12_335/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 31.235 74.695 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_335/VNB
  PIN sky130_ef_sc_hd__decap_12_334/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 31.235 80.215 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_334/VNB
  PIN sky130_ef_sc_hd__decap_12_333/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 31.235 85.735 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_333/VNB
  PIN sky130_fd_sc_hd__decap_6_53/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 31.235 91.255 31.405 ;
    END
  END sky130_fd_sc_hd__decap_6_53/VNB
  PIN sky130_fd_sc_hd__fill_1_101/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 31.265 93.960 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_101/VNB
  PIN sky130_ef_sc_hd__decap_12_332/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 31.235 94.935 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_332/VNB
  PIN sky130_ef_sc_hd__decap_12_331/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 31.235 100.455 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_331/VNB
  PIN sky130_ef_sc_hd__decap_12_330/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 31.235 105.975 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_330/VNB
  PIN sky130_ef_sc_hd__decap_12_329/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 31.235 111.495 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_329/VNB
  PIN sky130_fd_sc_hd__decap_6_52/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 31.235 117.015 31.405 ;
    END
  END sky130_fd_sc_hd__decap_6_52/VNB
  PIN sky130_fd_sc_hd__fill_1_100/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 31.265 119.720 31.375 ;
    END
  END sky130_fd_sc_hd__fill_1_100/VNB
  PIN sky130_ef_sc_hd__decap_12_328/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 31.235 120.695 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_328/VNB
  PIN sky130_ef_sc_hd__decap_12_327/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 31.235 126.215 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_327/VNB
  PIN sky130_ef_sc_hd__decap_12_326/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 31.235 131.735 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_326/VNB
  PIN sky130_ef_sc_hd__decap_12_325/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 31.235 137.255 31.405 ;
    END
  END sky130_ef_sc_hd__decap_12_325/VNB
  PIN sky130_ef_sc_hd__decap_12_324/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 36.675 57.215 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_324/VNB
  PIN sky130_fd_sc_hd__decap_3_54/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 36.675 55.835 36.845 ;
    END
  END sky130_fd_sc_hd__decap_3_54/VNB
  PIN sky130_ef_sc_hd__decap_12_323/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 36.675 62.735 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_323/VNB
  PIN sky130_ef_sc_hd__decap_12_322/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 36.815 68.255 36.845 ;
        RECT 68.080 36.705 68.255 36.815 ;
        RECT 68.085 36.675 68.255 36.705 ;
    END
  END sky130_ef_sc_hd__decap_12_322/VNB
  PIN sky130_ef_sc_hd__decap_12_321/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 36.675 73.775 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_321/VNB
  PIN sky130_fd_sc_hd__decap_4_9/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 36.675 79.295 36.845 ;
    END
  END sky130_fd_sc_hd__decap_4_9/VNB
  PIN sky130_fd_sc_hd__fill_1_98/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 36.705 81.080 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_98/VNB
  PIN sky130_ef_sc_hd__decap_12_320/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 36.675 82.055 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_320/VNB
  PIN sky130_ef_sc_hd__decap_12_319/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 36.675 87.575 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_319/VNB
  PIN sky130_ef_sc_hd__decap_12_318/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 36.675 93.095 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_318/VNB
  PIN sky130_ef_sc_hd__decap_12_317/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 36.675 98.615 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_317/VNB
  PIN sky130_fd_sc_hd__decap_6_51/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 36.675 104.135 36.845 ;
    END
  END sky130_fd_sc_hd__decap_6_51/VNB
  PIN sky130_fd_sc_hd__fill_1_97/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 36.705 106.840 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_97/VNB
  PIN sky130_ef_sc_hd__decap_12_316/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 36.675 107.815 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_316/VNB
  PIN sky130_ef_sc_hd__decap_12_315/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 36.675 113.335 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_315/VNB
  PIN sky130_ef_sc_hd__decap_12_314/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 36.675 118.855 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_314/VNB
  PIN sky130_ef_sc_hd__decap_12_313/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 36.675 124.375 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_313/VNB
  PIN sky130_fd_sc_hd__decap_6_50/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 36.675 129.895 36.845 ;
    END
  END sky130_fd_sc_hd__decap_6_50/VNB
  PIN sky130_fd_sc_hd__fill_1_96/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 36.705 132.600 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_96/VNB
  PIN sky130_ef_sc_hd__decap_12_312/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 36.675 133.575 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_312/VNB
  PIN sky130_fd_sc_hd__decap_8_17/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 36.675 139.095 36.845 ;
    END
  END sky130_fd_sc_hd__decap_8_17/VNB
  PIN sky130_fd_sc_hd__fill_1_95/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 36.705 142.720 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_95/VNB
  PIN sky130_fd_sc_hd__decap_3_53/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 36.675 144.155 36.845 ;
    END
  END sky130_fd_sc_hd__decap_3_53/VNB
  PIN sky130_ef_sc_hd__decap_12_309/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 36.675 69.175 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_309/VNB
  PIN sky130_ef_sc_hd__decap_12_308/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 36.675 74.695 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_308/VNB
  PIN sky130_ef_sc_hd__decap_12_307/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 36.675 80.215 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_307/VNB
  PIN sky130_ef_sc_hd__decap_12_306/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 36.675 85.735 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_306/VNB
  PIN sky130_fd_sc_hd__decap_6_49/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 36.675 91.255 36.845 ;
    END
  END sky130_fd_sc_hd__decap_6_49/VNB
  PIN sky130_fd_sc_hd__fill_1_93/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 36.705 93.960 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_93/VNB
  PIN sky130_ef_sc_hd__decap_12_305/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 36.675 94.935 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_305/VNB
  PIN sky130_ef_sc_hd__decap_12_304/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 36.675 100.455 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_304/VNB
  PIN sky130_ef_sc_hd__decap_12_303/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 36.675 105.975 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_303/VNB
  PIN sky130_ef_sc_hd__decap_12_302/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 36.675 111.495 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_302/VNB
  PIN sky130_fd_sc_hd__decap_6_48/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 36.675 117.015 36.845 ;
    END
  END sky130_fd_sc_hd__decap_6_48/VNB
  PIN sky130_fd_sc_hd__fill_1_92/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 36.705 119.720 36.815 ;
    END
  END sky130_fd_sc_hd__fill_1_92/VNB
  PIN sky130_ef_sc_hd__decap_12_301/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 36.675 120.695 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_301/VNB
  PIN sky130_ef_sc_hd__decap_12_300/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 36.675 126.215 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_300/VNB
  PIN sky130_ef_sc_hd__decap_12_299/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 36.675 131.735 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_299/VNB
  PIN sky130_ef_sc_hd__decap_12_298/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 36.675 137.255 36.845 ;
    END
  END sky130_ef_sc_hd__decap_12_298/VNB
  PIN sky130_ef_sc_hd__decap_12_297/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 42.115 57.215 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_297/VNB
  PIN sky130_fd_sc_hd__decap_3_50/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 42.115 55.835 42.285 ;
    END
  END sky130_fd_sc_hd__decap_3_50/VNB
  PIN sky130_ef_sc_hd__decap_12_296/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 42.115 62.735 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_296/VNB
  PIN sky130_ef_sc_hd__decap_12_295/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 42.255 68.255 42.285 ;
        RECT 68.080 42.145 68.255 42.255 ;
        RECT 68.085 42.115 68.255 42.145 ;
    END
  END sky130_ef_sc_hd__decap_12_295/VNB
  PIN sky130_ef_sc_hd__decap_12_294/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 42.115 73.775 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_294/VNB
  PIN sky130_fd_sc_hd__decap_4_8/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 42.115 79.295 42.285 ;
    END
  END sky130_fd_sc_hd__decap_4_8/VNB
  PIN sky130_fd_sc_hd__fill_1_90/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 42.145 81.080 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_90/VNB
  PIN sky130_ef_sc_hd__decap_12_293/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 42.115 82.055 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_293/VNB
  PIN sky130_ef_sc_hd__decap_12_292/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 42.115 87.575 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_292/VNB
  PIN sky130_ef_sc_hd__decap_12_291/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 42.115 93.095 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_291/VNB
  PIN sky130_ef_sc_hd__decap_12_290/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 42.115 98.615 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_290/VNB
  PIN sky130_fd_sc_hd__decap_6_47/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 42.115 104.135 42.285 ;
    END
  END sky130_fd_sc_hd__decap_6_47/VNB
  PIN sky130_fd_sc_hd__fill_1_89/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 42.145 106.840 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_89/VNB
  PIN sky130_ef_sc_hd__decap_12_289/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 42.115 107.815 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_289/VNB
  PIN sky130_ef_sc_hd__decap_12_288/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 42.115 113.335 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_288/VNB
  PIN sky130_ef_sc_hd__decap_12_287/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 42.115 118.855 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_287/VNB
  PIN sky130_ef_sc_hd__decap_12_286/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 42.115 124.375 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_286/VNB
  PIN sky130_fd_sc_hd__decap_6_46/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 42.115 129.895 42.285 ;
    END
  END sky130_fd_sc_hd__decap_6_46/VNB
  PIN sky130_fd_sc_hd__fill_1_88/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 42.145 132.600 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_88/VNB
  PIN sky130_ef_sc_hd__decap_12_285/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 42.115 133.575 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_285/VNB
  PIN sky130_fd_sc_hd__decap_8_16/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 42.115 139.095 42.285 ;
    END
  END sky130_fd_sc_hd__decap_8_16/VNB
  PIN sky130_fd_sc_hd__fill_1_87/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 42.145 142.720 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_87/VNB
  PIN sky130_fd_sc_hd__decap_3_49/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 42.115 144.155 42.285 ;
    END
  END sky130_fd_sc_hd__decap_3_49/VNB
  PIN sky130_ef_sc_hd__decap_12_283/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 47.555 57.215 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_283/VNB
  PIN sky130_fd_sc_hd__decap_3_47/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 47.555 55.835 47.725 ;
    END
  END sky130_fd_sc_hd__decap_3_47/VNB
  PIN sky130_ef_sc_hd__decap_12_281/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 47.555 62.735 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_281/VNB
  PIN sky130_ef_sc_hd__decap_12_280/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 42.115 69.175 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_280/VNB
  PIN sky130_ef_sc_hd__decap_12_279/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 47.695 68.255 47.725 ;
        RECT 68.080 47.585 68.255 47.695 ;
        RECT 68.085 47.555 68.255 47.585 ;
    END
  END sky130_ef_sc_hd__decap_12_279/VNB
  PIN sky130_ef_sc_hd__decap_12_278/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 42.115 74.695 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_278/VNB
  PIN sky130_ef_sc_hd__decap_12_277/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 47.555 73.775 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_277/VNB
  PIN sky130_fd_sc_hd__decap_4_7/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 47.555 79.295 47.725 ;
    END
  END sky130_fd_sc_hd__decap_4_7/VNB
  PIN sky130_ef_sc_hd__decap_12_276/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 42.115 80.215 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_276/VNB
  PIN sky130_fd_sc_hd__fill_1_85/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 47.585 81.080 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_85/VNB
  PIN sky130_ef_sc_hd__decap_12_275/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 47.555 82.055 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_275/VNB
  PIN sky130_ef_sc_hd__decap_12_274/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 42.115 85.735 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_274/VNB
  PIN sky130_fd_sc_hd__decap_6_45/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 42.115 91.255 42.285 ;
    END
  END sky130_fd_sc_hd__decap_6_45/VNB
  PIN sky130_ef_sc_hd__decap_12_273/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 47.555 87.575 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_273/VNB
  PIN sky130_fd_sc_hd__fill_1_84/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 42.145 93.960 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_84/VNB
  PIN sky130_ef_sc_hd__decap_12_272/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 42.115 94.935 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_272/VNB
  PIN sky130_ef_sc_hd__decap_12_271/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 47.555 93.095 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_271/VNB
  PIN sky130_ef_sc_hd__decap_12_270/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 42.115 100.455 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_270/VNB
  PIN sky130_ef_sc_hd__decap_12_269/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 47.555 98.615 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_269/VNB
  PIN sky130_ef_sc_hd__decap_12_268/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 42.115 105.975 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_268/VNB
  PIN sky130_fd_sc_hd__decap_6_44/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 47.555 104.135 47.725 ;
    END
  END sky130_fd_sc_hd__decap_6_44/VNB
  PIN sky130_fd_sc_hd__fill_1_83/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 47.585 106.840 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_83/VNB
  PIN sky130_ef_sc_hd__decap_12_267/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 47.555 107.815 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_267/VNB
  PIN sky130_ef_sc_hd__decap_12_266/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 42.115 111.495 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_266/VNB
  PIN sky130_ef_sc_hd__decap_12_265/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 47.555 113.335 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_265/VNB
  PIN sky130_fd_sc_hd__decap_6_43/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 42.115 117.015 42.285 ;
    END
  END sky130_fd_sc_hd__decap_6_43/VNB
  PIN sky130_fd_sc_hd__fill_1_82/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 42.145 119.720 42.255 ;
    END
  END sky130_fd_sc_hd__fill_1_82/VNB
  PIN sky130_ef_sc_hd__decap_12_264/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 42.115 120.695 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_264/VNB
  PIN sky130_ef_sc_hd__decap_12_263/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 47.555 118.855 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_263/VNB
  PIN sky130_ef_sc_hd__decap_12_262/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 42.115 126.215 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_262/VNB
  PIN sky130_ef_sc_hd__decap_12_261/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 47.555 124.375 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_261/VNB
  PIN sky130_ef_sc_hd__decap_12_260/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 42.115 131.735 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_260/VNB
  PIN sky130_fd_sc_hd__decap_6_42/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 47.555 129.895 47.725 ;
    END
  END sky130_fd_sc_hd__decap_6_42/VNB
  PIN sky130_ef_sc_hd__decap_12_259/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 42.115 137.255 42.285 ;
    END
  END sky130_ef_sc_hd__decap_12_259/VNB
  PIN sky130_fd_sc_hd__fill_1_81/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 47.585 132.600 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_81/VNB
  PIN sky130_ef_sc_hd__decap_12_258/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 47.555 133.575 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_258/VNB
  PIN sky130_fd_sc_hd__decap_8_15/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 47.555 139.095 47.725 ;
    END
  END sky130_fd_sc_hd__decap_8_15/VNB
  PIN sky130_fd_sc_hd__fill_1_79/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 47.585 142.720 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_79/VNB
  PIN sky130_fd_sc_hd__decap_3_45/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 47.555 144.155 47.725 ;
    END
  END sky130_fd_sc_hd__decap_3_45/VNB
  PIN sky130_ef_sc_hd__decap_12_255/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 47.555 69.175 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_255/VNB
  PIN sky130_ef_sc_hd__decap_12_254/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 47.555 74.695 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_254/VNB
  PIN sky130_ef_sc_hd__decap_12_253/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 47.555 80.215 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_253/VNB
  PIN sky130_ef_sc_hd__decap_12_252/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 47.555 85.735 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_252/VNB
  PIN sky130_fd_sc_hd__decap_6_41/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 47.555 91.255 47.725 ;
    END
  END sky130_fd_sc_hd__decap_6_41/VNB
  PIN sky130_fd_sc_hd__fill_1_77/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 47.585 93.960 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_77/VNB
  PIN sky130_ef_sc_hd__decap_12_251/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 47.555 94.935 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_251/VNB
  PIN sky130_ef_sc_hd__decap_12_250/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 47.555 100.455 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_250/VNB
  PIN sky130_ef_sc_hd__decap_12_249/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 47.555 105.975 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_249/VNB
  PIN sky130_ef_sc_hd__decap_12_248/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 47.555 111.495 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_248/VNB
  PIN sky130_fd_sc_hd__decap_6_40/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 47.555 117.015 47.725 ;
    END
  END sky130_fd_sc_hd__decap_6_40/VNB
  PIN sky130_fd_sc_hd__fill_1_76/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 47.585 119.720 47.695 ;
    END
  END sky130_fd_sc_hd__fill_1_76/VNB
  PIN sky130_ef_sc_hd__decap_12_247/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 47.555 120.695 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_247/VNB
  PIN sky130_ef_sc_hd__decap_12_246/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 47.555 126.215 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_246/VNB
  PIN sky130_ef_sc_hd__decap_12_245/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 47.555 131.735 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_245/VNB
  PIN sky130_ef_sc_hd__decap_12_244/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 47.555 137.255 47.725 ;
    END
  END sky130_ef_sc_hd__decap_12_244/VNB
  PIN sky130_ef_sc_hd__decap_12_243/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 52.995 57.215 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_243/VNB
  PIN sky130_fd_sc_hd__decap_3_42/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 52.995 55.835 53.165 ;
    END
  END sky130_fd_sc_hd__decap_3_42/VNB
  PIN sky130_ef_sc_hd__decap_12_242/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 52.995 62.735 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_242/VNB
  PIN sky130_ef_sc_hd__decap_12_241/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 53.135 68.255 53.165 ;
        RECT 68.080 53.025 68.255 53.135 ;
        RECT 68.085 52.995 68.255 53.025 ;
    END
  END sky130_ef_sc_hd__decap_12_241/VNB
  PIN sky130_ef_sc_hd__decap_12_240/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 52.995 73.775 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_240/VNB
  PIN sky130_fd_sc_hd__decap_4_6/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 52.995 79.295 53.165 ;
    END
  END sky130_fd_sc_hd__decap_4_6/VNB
  PIN sky130_fd_sc_hd__fill_1_74/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 53.025 81.080 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_74/VNB
  PIN sky130_ef_sc_hd__decap_12_239/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 52.995 82.055 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_239/VNB
  PIN sky130_ef_sc_hd__decap_12_238/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 52.995 87.575 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_238/VNB
  PIN sky130_ef_sc_hd__decap_12_237/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 52.995 93.095 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_237/VNB
  PIN sky130_ef_sc_hd__decap_12_236/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 52.995 98.615 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_236/VNB
  PIN sky130_fd_sc_hd__decap_6_39/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 52.995 104.135 53.165 ;
    END
  END sky130_fd_sc_hd__decap_6_39/VNB
  PIN sky130_fd_sc_hd__fill_1_73/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 53.025 106.840 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_73/VNB
  PIN sky130_ef_sc_hd__decap_12_235/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 52.995 107.815 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_235/VNB
  PIN sky130_ef_sc_hd__decap_12_234/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 52.995 113.335 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_234/VNB
  PIN sky130_ef_sc_hd__decap_12_233/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 52.995 118.855 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_233/VNB
  PIN sky130_ef_sc_hd__decap_12_232/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 52.995 124.375 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_232/VNB
  PIN sky130_fd_sc_hd__decap_6_38/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 52.995 129.895 53.165 ;
    END
  END sky130_fd_sc_hd__decap_6_38/VNB
  PIN sky130_fd_sc_hd__fill_1_72/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 53.025 132.600 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_72/VNB
  PIN sky130_ef_sc_hd__decap_12_231/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 52.995 133.575 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_231/VNB
  PIN sky130_fd_sc_hd__decap_8_14/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 52.995 139.095 53.165 ;
    END
  END sky130_fd_sc_hd__decap_8_14/VNB
  PIN sky130_fd_sc_hd__fill_1_71/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 53.025 142.720 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_71/VNB
  PIN sky130_fd_sc_hd__decap_3_41/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 52.995 144.155 53.165 ;
    END
  END sky130_fd_sc_hd__decap_3_41/VNB
  PIN sky130_fd_sc_hd__buf_1_2/X
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 66.205 54.640 66.475 55.545 ;
        RECT 66.295 53.840 66.475 54.640 ;
        RECT 66.215 53.335 66.475 53.840 ;
    END
  END sky130_fd_sc_hd__buf_1_2/X
  PIN sky130_fd_sc_hd__buf_1_2/A
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 65.295 57.695 65.550 58.265 ;
        RECT 65.380 57.025 65.550 57.695 ;
        RECT 65.215 56.055 65.550 57.025 ;
        RECT 65.285 54.065 65.625 54.435 ;
      LAYER mcon ;
        RECT 65.325 56.225 65.495 56.395 ;
        RECT 65.325 54.185 65.495 54.355 ;
      LAYER met1 ;
        RECT 65.250 56.180 65.570 56.440 ;
        RECT 65.250 54.140 65.570 54.400 ;
      LAYER via ;
        RECT 65.280 56.180 65.540 56.440 ;
        RECT 65.280 54.140 65.540 54.400 ;
      LAYER met2 ;
        RECT 65.280 56.150 65.540 56.470 ;
        RECT 65.340 54.430 65.480 56.150 ;
        RECT 65.280 54.110 65.540 54.430 ;
    END
  END sky130_fd_sc_hd__buf_1_2/A
  PIN sky130_fd_sc_hd__buf_1_2/VNB
    PORT
      LAYER pwell ;
        RECT 65.335 52.995 65.505 53.165 ;
    END
  END sky130_fd_sc_hd__buf_1_2/VNB
  PIN sky130_fd_sc_hd__inv_2_4/A
    ANTENNAGATEAREA 0.868500 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 57.925 65.520 58.195 66.425 ;
        RECT 58.015 64.720 58.195 65.520 ;
        RECT 57.935 64.215 58.195 64.720 ;
        RECT 66.665 59.595 67.000 59.845 ;
        RECT 63.375 58.095 63.650 58.265 ;
        RECT 63.375 57.925 63.655 58.095 ;
        RECT 63.375 57.105 63.650 57.925 ;
        RECT 66.665 54.155 66.995 54.405 ;
      LAYER mcon ;
        RECT 57.965 64.385 58.135 64.555 ;
        RECT 66.705 59.625 66.875 59.795 ;
        RECT 63.485 57.925 63.655 58.095 ;
        RECT 66.705 54.185 66.875 54.355 ;
      LAYER met1 ;
        RECT 57.905 64.540 58.195 64.585 ;
        RECT 63.410 64.540 63.730 64.600 ;
        RECT 57.905 64.400 63.730 64.540 ;
        RECT 57.905 64.355 58.195 64.400 ;
        RECT 63.410 64.340 63.730 64.400 ;
        RECT 63.410 59.780 63.730 59.840 ;
        RECT 66.645 59.780 66.935 59.825 ;
        RECT 63.410 59.640 66.935 59.780 ;
        RECT 63.410 59.580 63.730 59.640 ;
        RECT 66.645 59.595 66.935 59.640 ;
        RECT 63.410 57.880 63.730 58.140 ;
        RECT 63.870 54.680 64.190 54.740 ;
        RECT 63.870 54.540 66.860 54.680 ;
        RECT 63.870 54.480 64.190 54.540 ;
        RECT 66.720 54.385 66.860 54.540 ;
        RECT 66.645 54.155 66.935 54.385 ;
      LAYER via ;
        RECT 63.440 64.340 63.700 64.600 ;
        RECT 63.440 59.580 63.700 59.840 ;
        RECT 63.440 57.880 63.700 58.140 ;
        RECT 63.900 54.480 64.160 54.740 ;
      LAYER met2 ;
        RECT 63.440 64.310 63.700 64.630 ;
        RECT 63.500 59.870 63.640 64.310 ;
        RECT 63.440 59.550 63.700 59.870 ;
        RECT 63.500 58.170 63.640 59.550 ;
        RECT 63.440 57.850 63.700 58.170 ;
        RECT 63.500 56.890 63.640 57.850 ;
        RECT 63.500 56.750 64.100 56.890 ;
        RECT 63.960 54.770 64.100 56.750 ;
        RECT 63.900 54.450 64.160 54.770 ;
    END
  END sky130_fd_sc_hd__inv_2_4/A
  PIN sky130_fd_sc_hd__inv_2_4/Y
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 67.630 57.415 67.905 58.265 ;
        RECT 67.625 57.245 67.905 57.415 ;
        RECT 67.630 57.105 67.905 57.245 ;
        RECT 67.085 54.565 67.415 55.545 ;
        RECT 67.165 53.965 67.415 54.565 ;
        RECT 67.085 53.335 67.415 53.965 ;
      LAYER mcon ;
        RECT 67.165 55.205 67.335 55.375 ;
      LAYER met1 ;
        RECT 67.550 57.200 67.870 57.460 ;
        RECT 67.105 55.360 67.395 55.405 ;
        RECT 67.550 55.360 67.870 55.420 ;
        RECT 67.105 55.220 67.870 55.360 ;
        RECT 67.105 55.175 67.395 55.220 ;
        RECT 67.550 55.160 67.870 55.220 ;
      LAYER via ;
        RECT 67.580 57.200 67.840 57.460 ;
        RECT 67.580 55.160 67.840 55.420 ;
      LAYER met2 ;
        RECT 67.580 57.170 67.840 57.490 ;
        RECT 67.640 55.450 67.780 57.170 ;
        RECT 67.580 55.130 67.840 55.450 ;
    END
  END sky130_fd_sc_hd__inv_2_4/Y
  PIN sky130_fd_sc_hd__inv_2_4/VNB
    PORT
      LAYER pwell ;
        RECT 66.705 52.995 66.875 53.165 ;
    END
  END sky130_fd_sc_hd__inv_2_4/VNB
  PIN sky130_ef_sc_hd__decap_12_229/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 52.995 69.175 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_229/VNB
  PIN sky130_ef_sc_hd__decap_12_228/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 52.995 74.695 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_228/VNB
  PIN sky130_ef_sc_hd__decap_12_227/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 52.995 80.215 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_227/VNB
  PIN sky130_ef_sc_hd__decap_12_226/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 52.995 85.735 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_226/VNB
  PIN sky130_fd_sc_hd__decap_6_36/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 52.995 91.255 53.165 ;
    END
  END sky130_fd_sc_hd__decap_6_36/VNB
  PIN sky130_fd_sc_hd__fill_1_69/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 53.025 93.960 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_69/VNB
  PIN sky130_ef_sc_hd__decap_12_225/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 52.995 94.935 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_225/VNB
  PIN sky130_ef_sc_hd__decap_12_224/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 52.995 100.455 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_224/VNB
  PIN sky130_ef_sc_hd__decap_12_223/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 52.995 105.975 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_223/VNB
  PIN sky130_ef_sc_hd__decap_12_222/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 52.995 111.495 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_222/VNB
  PIN sky130_fd_sc_hd__decap_6_35/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 52.995 117.015 53.165 ;
    END
  END sky130_fd_sc_hd__decap_6_35/VNB
  PIN sky130_fd_sc_hd__fill_1_68/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 53.025 119.720 53.135 ;
    END
  END sky130_fd_sc_hd__fill_1_68/VNB
  PIN sky130_ef_sc_hd__decap_12_221/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 52.995 120.695 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_221/VNB
  PIN sky130_ef_sc_hd__decap_12_220/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 52.995 126.215 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_220/VNB
  PIN sky130_ef_sc_hd__decap_12_219/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 52.995 131.735 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_219/VNB
  PIN sky130_ef_sc_hd__decap_12_218/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 52.995 137.255 53.165 ;
    END
  END sky130_ef_sc_hd__decap_12_218/VNB
  PIN sky130_fd_sc_hd__decap_8_13/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 58.435 57.215 58.605 ;
    END
  END sky130_fd_sc_hd__decap_8_13/VNB
  PIN sky130_fd_sc_hd__decap_3_38/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 58.435 55.835 58.605 ;
    END
  END sky130_fd_sc_hd__decap_3_38/VNB
  PIN sky130_fd_sc_hd__fill_2_4/VNB
    PORT
      LAYER pwell ;
        RECT 60.735 58.460 60.895 58.570 ;
    END
  END sky130_fd_sc_hd__fill_2_4/VNB
  PIN sky130_fd_sc_hd__mux2_1_0/S
    ANTENNAGATEAREA 1.440000 ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER li1 ;
        RECT 66.075 68.495 66.935 68.745 ;
        RECT 66.655 67.905 66.935 68.495 ;
        RECT 67.970 68.125 68.300 68.635 ;
        RECT 65.235 67.735 66.935 67.905 ;
        RECT 65.235 66.935 65.565 67.735 ;
        RECT 66.075 66.935 66.405 67.735 ;
        RECT 64.535 57.195 64.730 57.525 ;
        RECT 66.550 57.195 66.745 57.525 ;
        RECT 69.885 57.195 70.215 57.445 ;
        RECT 62.095 56.890 62.845 57.080 ;
        RECT 62.675 56.225 62.845 56.890 ;
        RECT 64.535 56.225 64.705 57.195 ;
        RECT 62.675 56.055 64.705 56.225 ;
        RECT 66.575 56.225 66.745 57.195 ;
        RECT 68.435 56.890 69.185 57.080 ;
        RECT 68.435 56.225 68.605 56.890 ;
        RECT 66.575 56.055 68.605 56.225 ;
      LAYER mcon ;
        RECT 66.705 68.465 66.875 68.635 ;
        RECT 68.085 68.465 68.255 68.635 ;
        RECT 69.925 57.245 70.095 57.415 ;
        RECT 62.565 56.905 62.735 57.075 ;
        RECT 68.545 56.905 68.715 57.075 ;
      LAYER met1 ;
        RECT 66.645 68.620 66.935 68.665 ;
        RECT 68.025 68.620 68.315 68.665 ;
        RECT 68.470 68.620 68.790 68.680 ;
        RECT 66.645 68.480 68.790 68.620 ;
        RECT 66.645 68.435 66.935 68.480 ;
        RECT 68.025 68.435 68.315 68.480 ;
        RECT 68.470 68.420 68.790 68.480 ;
        RECT 69.865 57.400 70.155 57.445 ;
        RECT 68.560 57.260 70.155 57.400 ;
        RECT 68.560 57.120 68.700 57.260 ;
        RECT 69.865 57.215 70.155 57.260 ;
        RECT 62.505 57.060 62.795 57.105 ;
        RECT 68.470 57.060 68.790 57.120 ;
        RECT 62.505 56.920 68.790 57.060 ;
        RECT 62.505 56.875 62.795 56.920 ;
        RECT 68.470 56.860 68.790 56.920 ;
      LAYER via ;
        RECT 68.500 68.420 68.760 68.680 ;
        RECT 68.500 56.860 68.760 57.120 ;
      LAYER met2 ;
        RECT 68.500 68.390 68.760 68.710 ;
        RECT 68.560 57.150 68.700 68.390 ;
        RECT 68.500 56.830 68.760 57.150 ;
    END
  END sky130_fd_sc_hd__mux2_1_0/S
  PIN sky130_fd_sc_hd__mux2_1_0/A1
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 67.075 60.005 67.405 60.985 ;
        RECT 67.170 59.405 67.340 60.005 ;
        RECT 66.645 58.775 67.340 59.405 ;
        RECT 63.015 56.905 63.205 58.265 ;
        RECT 63.855 56.905 64.025 57.705 ;
        RECT 71.265 57.195 71.595 57.445 ;
        RECT 63.015 56.735 64.025 56.905 ;
      LAYER mcon ;
        RECT 66.705 58.945 66.875 59.115 ;
        RECT 63.025 57.925 63.195 58.095 ;
        RECT 71.305 57.245 71.475 57.415 ;
      LAYER met1 ;
        RECT 62.950 59.100 63.270 59.160 ;
        RECT 66.645 59.100 66.935 59.145 ;
        RECT 71.230 59.100 71.550 59.160 ;
        RECT 62.950 58.960 71.550 59.100 ;
        RECT 62.950 58.900 63.270 58.960 ;
        RECT 66.645 58.915 66.935 58.960 ;
        RECT 71.230 58.900 71.550 58.960 ;
        RECT 62.950 57.880 63.270 58.140 ;
        RECT 71.230 57.200 71.550 57.460 ;
      LAYER via ;
        RECT 62.980 58.900 63.240 59.160 ;
        RECT 71.260 58.900 71.520 59.160 ;
        RECT 62.980 57.880 63.240 58.140 ;
        RECT 71.260 57.200 71.520 57.460 ;
      LAYER met2 ;
        RECT 62.980 58.870 63.240 59.190 ;
        RECT 71.260 58.870 71.520 59.190 ;
        RECT 63.040 58.170 63.180 58.870 ;
        RECT 62.980 57.850 63.240 58.170 ;
        RECT 71.320 57.490 71.460 58.870 ;
        RECT 71.260 57.170 71.520 57.490 ;
    END
  END sky130_fd_sc_hd__mux2_1_0/A1
  PIN sky130_fd_sc_hd__mux2_1_0/VNB
    PORT
      LAYER pwell ;
        RECT 65.050 58.435 65.220 58.605 ;
    END
  END sky130_fd_sc_hd__mux2_1_0/VNB
  PIN sky130_fd_sc_hd__mux2_1_1/A1
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 67.255 56.905 67.425 57.705 ;
        RECT 68.075 56.905 68.265 58.265 ;
        RECT 71.685 57.635 72.015 58.265 ;
        RECT 71.765 57.035 72.015 57.635 ;
        RECT 67.255 56.735 68.265 56.905 ;
        RECT 71.685 56.055 72.015 57.035 ;
      LAYER mcon ;
        RECT 68.085 57.585 68.255 57.755 ;
        RECT 71.765 57.585 71.935 57.755 ;
      LAYER met1 ;
        RECT 68.025 57.740 68.315 57.785 ;
        RECT 71.705 57.740 71.995 57.785 ;
        RECT 68.025 57.600 71.995 57.740 ;
        RECT 68.025 57.555 68.315 57.600 ;
        RECT 71.705 57.555 71.995 57.600 ;
    END
  END sky130_fd_sc_hd__mux2_1_1/A1
  PIN sky130_fd_sc_hd__mux2_1_1/X
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 65.745 62.605 66.075 62.975 ;
        RECT 65.730 57.695 65.985 58.265 ;
        RECT 65.730 57.025 65.900 57.695 ;
        RECT 65.730 56.055 66.065 57.025 ;
      LAYER mcon ;
        RECT 65.785 62.685 65.955 62.855 ;
        RECT 65.785 57.925 65.955 58.095 ;
      LAYER met1 ;
        RECT 65.250 62.840 65.570 62.900 ;
        RECT 65.725 62.840 66.015 62.885 ;
        RECT 65.250 62.700 66.015 62.840 ;
        RECT 65.250 62.640 65.570 62.700 ;
        RECT 65.725 62.655 66.015 62.700 ;
        RECT 65.250 58.080 65.570 58.140 ;
        RECT 65.725 58.080 66.015 58.125 ;
        RECT 65.250 57.940 66.015 58.080 ;
        RECT 65.250 57.880 65.570 57.940 ;
        RECT 65.725 57.895 66.015 57.940 ;
      LAYER via ;
        RECT 65.280 62.640 65.540 62.900 ;
        RECT 65.280 57.880 65.540 58.140 ;
      LAYER met2 ;
        RECT 65.280 62.610 65.540 62.930 ;
        RECT 65.340 58.170 65.480 62.610 ;
        RECT 65.280 57.850 65.540 58.170 ;
    END
  END sky130_fd_sc_hd__mux2_1_1/X
  PIN sky130_fd_sc_hd__mux2_1_1/VNB
    PORT
      LAYER pwell ;
        RECT 66.060 58.435 66.230 58.605 ;
    END
  END sky130_fd_sc_hd__mux2_1_1/VNB
  PIN sky130_fd_sc_hd__inv_2_3/Y
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 70.305 57.635 70.635 58.265 ;
        RECT 70.385 57.035 70.635 57.635 ;
        RECT 70.305 56.055 70.635 57.035 ;
    END
  END sky130_fd_sc_hd__inv_2_3/Y
  PIN sky130_fd_sc_hd__inv_2_3/VNB
    PORT
      LAYER pwell ;
        RECT 69.925 58.435 70.095 58.605 ;
    END
  END sky130_fd_sc_hd__inv_2_3/VNB
  PIN sky130_fd_sc_hd__inv_2_2/VNB
    PORT
      LAYER pwell ;
        RECT 71.305 58.435 71.475 58.605 ;
    END
  END sky130_fd_sc_hd__inv_2_2/VNB
  PIN sky130_ef_sc_hd__decap_12_217/VNB
    PORT
      LAYER pwell ;
        RECT 72.685 58.435 72.855 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_217/VNB
  PIN sky130_fd_sc_hd__decap_6_34/VNB
    PORT
      LAYER pwell ;
        RECT 78.205 58.435 78.375 58.605 ;
    END
  END sky130_fd_sc_hd__decap_6_34/VNB
  PIN sky130_fd_sc_hd__fill_1_66/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 58.465 81.080 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_66/VNB
  PIN sky130_ef_sc_hd__decap_12_216/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 58.435 82.055 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_216/VNB
  PIN sky130_ef_sc_hd__decap_12_215/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 58.435 87.575 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_215/VNB
  PIN sky130_ef_sc_hd__decap_12_214/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 58.435 93.095 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_214/VNB
  PIN sky130_ef_sc_hd__decap_12_213/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 58.435 98.615 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_213/VNB
  PIN sky130_fd_sc_hd__decap_6_33/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 58.435 104.135 58.605 ;
    END
  END sky130_fd_sc_hd__decap_6_33/VNB
  PIN sky130_fd_sc_hd__fill_1_65/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 58.465 106.840 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_65/VNB
  PIN sky130_ef_sc_hd__decap_12_212/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 58.435 107.815 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_212/VNB
  PIN sky130_ef_sc_hd__decap_12_211/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 58.435 113.335 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_211/VNB
  PIN sky130_ef_sc_hd__decap_12_210/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 58.435 118.855 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_210/VNB
  PIN sky130_ef_sc_hd__decap_12_209/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 58.435 124.375 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_209/VNB
  PIN sky130_fd_sc_hd__decap_6_32/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 58.435 129.895 58.605 ;
    END
  END sky130_fd_sc_hd__decap_6_32/VNB
  PIN sky130_fd_sc_hd__fill_1_64/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 58.465 132.600 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_64/VNB
  PIN sky130_ef_sc_hd__decap_12_208/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 58.435 133.575 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_208/VNB
  PIN sky130_fd_sc_hd__decap_8_12/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 58.435 139.095 58.605 ;
    END
  END sky130_fd_sc_hd__decap_8_12/VNB
  PIN sky130_fd_sc_hd__fill_1_63/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 58.465 142.720 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_63/VNB
  PIN sky130_fd_sc_hd__decap_3_37/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 58.435 144.155 58.605 ;
    END
  END sky130_fd_sc_hd__decap_3_37/VNB
  PIN sky130_fd_sc_hd__decap_8_11/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 58.435 62.735 58.605 ;
    END
  END sky130_fd_sc_hd__decap_8_11/VNB
  PIN sky130_fd_sc_hd__fill_1_62/VNB
    PORT
      LAYER pwell ;
        RECT 66.240 58.465 66.360 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_62/VNB
  PIN sky130_fd_sc_hd__nand2_1_1/B
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 70.345 73.515 70.675 73.765 ;
        RECT 63.360 70.475 63.695 70.725 ;
        RECT 70.315 68.545 71.075 68.765 ;
        RECT 65.735 68.075 66.485 68.325 ;
        RECT 70.845 67.955 71.075 68.545 ;
        RECT 68.925 67.775 71.075 67.955 ;
        RECT 68.925 67.635 70.645 67.775 ;
        RECT 70.315 67.275 70.645 67.635 ;
        RECT 67.510 59.575 67.845 59.845 ;
      LAYER mcon ;
        RECT 70.385 73.565 70.555 73.735 ;
        RECT 63.485 70.505 63.655 70.675 ;
        RECT 66.245 68.125 66.415 68.295 ;
        RECT 69.005 67.785 69.175 67.955 ;
        RECT 67.625 59.625 67.795 59.795 ;
      LAYER met1 ;
        RECT 68.930 73.720 69.250 73.780 ;
        RECT 70.325 73.720 70.615 73.765 ;
        RECT 68.930 73.580 70.615 73.720 ;
        RECT 68.930 73.520 69.250 73.580 ;
        RECT 70.325 73.535 70.615 73.580 ;
        RECT 63.425 70.660 63.715 70.705 ;
        RECT 65.250 70.660 65.570 70.720 ;
        RECT 63.425 70.520 65.570 70.660 ;
        RECT 63.425 70.475 63.715 70.520 ;
        RECT 65.250 70.460 65.570 70.520 ;
        RECT 65.250 68.280 65.570 68.340 ;
        RECT 66.185 68.280 66.475 68.325 ;
        RECT 65.250 68.140 66.475 68.280 ;
        RECT 65.250 68.080 65.570 68.140 ;
        RECT 66.185 68.095 66.475 68.140 ;
        RECT 66.260 67.600 66.400 68.095 ;
        RECT 68.930 67.740 69.250 68.000 ;
        RECT 69.020 67.600 69.160 67.740 ;
        RECT 66.260 67.460 69.160 67.600 ;
        RECT 67.565 59.780 67.855 59.825 ;
        RECT 68.930 59.780 69.250 59.840 ;
        RECT 67.565 59.640 69.250 59.780 ;
        RECT 67.565 59.595 67.855 59.640 ;
        RECT 68.930 59.580 69.250 59.640 ;
      LAYER via ;
        RECT 68.960 73.520 69.220 73.780 ;
        RECT 65.280 70.460 65.540 70.720 ;
        RECT 65.280 68.080 65.540 68.340 ;
        RECT 68.960 67.740 69.220 68.000 ;
        RECT 68.960 59.580 69.220 59.840 ;
      LAYER met2 ;
        RECT 68.960 73.490 69.220 73.810 ;
        RECT 65.280 70.430 65.540 70.750 ;
        RECT 65.340 68.370 65.480 70.430 ;
        RECT 65.280 68.050 65.540 68.370 ;
        RECT 69.020 68.030 69.160 73.490 ;
        RECT 68.960 67.710 69.220 68.030 ;
        RECT 69.020 59.870 69.160 67.710 ;
        RECT 68.960 59.550 69.220 59.870 ;
    END
  END sky130_fd_sc_hd__nand2_1_1/B
  PIN sky130_fd_sc_hd__nand2_1_1/VNB
    PORT
      LAYER pwell ;
        RECT 67.630 58.435 67.800 58.605 ;
    END
  END sky130_fd_sc_hd__nand2_1_1/VNB
  PIN sky130_fd_sc_hd__fill_1_61/VNB
    PORT
      LAYER pwell ;
        RECT 68.080 58.465 68.200 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_61/VNB
  PIN sky130_ef_sc_hd__decap_12_206/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 58.435 69.175 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_206/VNB
  PIN sky130_ef_sc_hd__decap_12_205/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 58.435 74.695 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_205/VNB
  PIN sky130_ef_sc_hd__decap_12_204/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 58.435 80.215 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_204/VNB
  PIN sky130_ef_sc_hd__decap_12_203/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 58.435 85.735 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_203/VNB
  PIN sky130_fd_sc_hd__decap_6_31/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 58.435 91.255 58.605 ;
    END
  END sky130_fd_sc_hd__decap_6_31/VNB
  PIN sky130_fd_sc_hd__fill_1_60/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 58.465 93.960 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_60/VNB
  PIN sky130_ef_sc_hd__decap_12_202/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 58.435 94.935 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_202/VNB
  PIN sky130_ef_sc_hd__decap_12_201/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 58.435 100.455 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_201/VNB
  PIN sky130_ef_sc_hd__decap_12_200/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 58.435 105.975 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_200/VNB
  PIN sky130_ef_sc_hd__decap_12_199/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 58.435 111.495 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_199/VNB
  PIN sky130_fd_sc_hd__decap_6_30/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 58.435 117.015 58.605 ;
    END
  END sky130_fd_sc_hd__decap_6_30/VNB
  PIN sky130_fd_sc_hd__fill_1_59/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 58.465 119.720 58.575 ;
    END
  END sky130_fd_sc_hd__fill_1_59/VNB
  PIN sky130_ef_sc_hd__decap_12_198/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 58.435 120.695 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_198/VNB
  PIN sky130_ef_sc_hd__decap_12_197/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 58.435 126.215 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_197/VNB
  PIN sky130_ef_sc_hd__decap_12_196/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 58.435 131.735 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_196/VNB
  PIN sky130_ef_sc_hd__decap_12_195/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 58.435 137.255 58.605 ;
    END
  END sky130_ef_sc_hd__decap_12_195/VNB
  PIN sky130_ef_sc_hd__decap_12_194/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 63.875 57.225 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_194/VNB
  PIN sky130_fd_sc_hd__decap_3_34/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 63.875 55.835 64.045 ;
    END
  END sky130_fd_sc_hd__decap_3_34/VNB
  PIN sky130_ef_sc_hd__decap_12_193/VNB
    PORT
      LAYER pwell ;
        RECT 58.425 63.875 58.595 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_193/VNB
  PIN sky130_fd_sc_hd__decap_6_29/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 63.875 62.735 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_29/VNB
  PIN sky130_fd_sc_hd__fill_1_57/VNB
    PORT
      LAYER pwell ;
        RECT 65.320 63.905 65.440 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_57/VNB
  PIN sky130_fd_sc_hd__clkbuf_1_0/X
    ANTENNAGATEAREA 0.318000 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 67.125 70.395 67.395 71.015 ;
        RECT 67.510 67.725 67.800 68.635 ;
        RECT 66.675 63.200 66.935 63.705 ;
        RECT 66.765 62.400 66.935 63.200 ;
        RECT 66.665 61.495 66.935 62.400 ;
      LAYER mcon ;
        RECT 67.165 70.505 67.335 70.675 ;
        RECT 67.625 67.785 67.795 67.955 ;
        RECT 66.705 63.365 66.875 63.535 ;
      LAYER met1 ;
        RECT 67.105 70.660 67.395 70.705 ;
        RECT 67.550 70.660 67.870 70.720 ;
        RECT 67.105 70.520 67.870 70.660 ;
        RECT 67.105 70.475 67.395 70.520 ;
        RECT 67.550 70.460 67.870 70.520 ;
        RECT 67.550 67.740 67.870 68.000 ;
        RECT 66.645 63.520 66.935 63.565 ;
        RECT 67.550 63.520 67.870 63.580 ;
        RECT 66.645 63.380 67.870 63.520 ;
        RECT 66.645 63.335 66.935 63.380 ;
        RECT 67.550 63.320 67.870 63.380 ;
      LAYER via ;
        RECT 67.580 70.460 67.840 70.720 ;
        RECT 67.580 67.740 67.840 68.000 ;
        RECT 67.580 63.320 67.840 63.580 ;
      LAYER met2 ;
        RECT 67.580 70.430 67.840 70.750 ;
        RECT 67.640 68.030 67.780 70.430 ;
        RECT 67.580 67.710 67.840 68.030 ;
        RECT 67.640 63.610 67.780 67.710 ;
        RECT 67.580 63.290 67.840 63.610 ;
    END
  END sky130_fd_sc_hd__clkbuf_1_0/X
  PIN sky130_fd_sc_hd__clkbuf_1_0/VNB
    PORT
      LAYER pwell ;
        RECT 65.785 63.875 65.955 64.045 ;
    END
  END sky130_fd_sc_hd__clkbuf_1_0/VNB
  PIN sky130_fd_sc_hd__decap_8_10/VNB
    PORT
      LAYER pwell ;
        RECT 63.945 63.875 64.115 64.045 ;
    END
  END sky130_fd_sc_hd__decap_8_10/VNB
  PIN sky130_ef_sc_hd__decap_12_192/VNB
    PORT
      LAYER pwell ;
        RECT 67.165 63.875 67.335 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_192/VNB
  PIN sky130_fd_sc_hd__fill_2_3/VNB
    PORT
      LAYER pwell ;
        RECT 67.635 63.910 67.795 64.020 ;
    END
  END sky130_fd_sc_hd__fill_2_3/VNB
  PIN sky130_ef_sc_hd__decap_12_190/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 63.875 69.175 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_190/VNB
  PIN sky130_ef_sc_hd__decap_12_191/VNB
    PORT
      LAYER pwell ;
        RECT 72.685 63.875 72.855 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_191/VNB
  PIN sky130_ef_sc_hd__decap_12_189/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 63.875 74.695 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_189/VNB
  PIN sky130_fd_sc_hd__decap_6_28/VNB
    PORT
      LAYER pwell ;
        RECT 78.205 63.875 78.375 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_28/VNB
  PIN sky130_fd_sc_hd__fill_1_56/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 63.905 81.080 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_56/VNB
  PIN sky130_ef_sc_hd__decap_12_188/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 63.875 82.055 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_188/VNB
  PIN sky130_ef_sc_hd__decap_12_187/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 63.875 80.215 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_187/VNB
  PIN sky130_ef_sc_hd__decap_12_186/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 63.875 87.575 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_186/VNB
  PIN sky130_ef_sc_hd__decap_12_185/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 63.875 85.735 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_185/VNB
  PIN sky130_fd_sc_hd__decap_6_27/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 63.875 91.255 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_27/VNB
  PIN sky130_fd_sc_hd__fill_1_55/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 63.905 93.960 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_55/VNB
  PIN sky130_ef_sc_hd__decap_12_184/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 63.875 93.095 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_184/VNB
  PIN sky130_ef_sc_hd__decap_12_183/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 63.875 94.935 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_183/VNB
  PIN sky130_ef_sc_hd__decap_12_182/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 63.875 98.615 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_182/VNB
  PIN sky130_ef_sc_hd__decap_12_181/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 63.875 100.455 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_181/VNB
  PIN sky130_fd_sc_hd__decap_6_26/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 63.875 104.135 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_26/VNB
  PIN sky130_fd_sc_hd__fill_1_54/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 63.905 106.840 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_54/VNB
  PIN sky130_ef_sc_hd__decap_12_180/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 63.875 107.815 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_180/VNB
  PIN sky130_ef_sc_hd__decap_12_179/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 63.875 105.975 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_179/VNB
  PIN sky130_ef_sc_hd__decap_12_178/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 63.875 113.335 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_178/VNB
  PIN sky130_ef_sc_hd__decap_12_177/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 63.875 111.495 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_177/VNB
  PIN sky130_ef_sc_hd__decap_12_176/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 63.875 118.855 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_176/VNB
  PIN sky130_fd_sc_hd__decap_6_25/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 63.875 117.015 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_25/VNB
  PIN sky130_fd_sc_hd__fill_1_53/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 63.905 119.720 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_53/VNB
  PIN sky130_ef_sc_hd__decap_12_175/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 63.875 120.695 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_175/VNB
  PIN sky130_ef_sc_hd__decap_12_174/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 63.875 124.375 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_174/VNB
  PIN sky130_ef_sc_hd__decap_12_173/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 63.875 126.215 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_173/VNB
  PIN sky130_fd_sc_hd__decap_6_24/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 63.875 129.895 64.045 ;
    END
  END sky130_fd_sc_hd__decap_6_24/VNB
  PIN sky130_ef_sc_hd__decap_12_172/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 63.875 131.735 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_172/VNB
  PIN sky130_fd_sc_hd__fill_1_52/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 63.905 132.600 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_52/VNB
  PIN sky130_ef_sc_hd__decap_12_171/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 63.875 133.575 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_171/VNB
  PIN sky130_ef_sc_hd__decap_12_170/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 63.875 137.255 64.045 ;
    END
  END sky130_ef_sc_hd__decap_12_170/VNB
  PIN sky130_fd_sc_hd__decap_8_9/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 63.875 139.095 64.045 ;
    END
  END sky130_fd_sc_hd__decap_8_9/VNB
  PIN sky130_fd_sc_hd__fill_1_51/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 63.905 142.720 64.015 ;
    END
  END sky130_fd_sc_hd__fill_1_51/VNB
  PIN sky130_fd_sc_hd__decap_3_32/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 63.875 144.155 64.045 ;
    END
  END sky130_fd_sc_hd__decap_3_32/VNB
  PIN sky130_ef_sc_hd__decap_12_169/VNB
    PORT
      LAYER pwell ;
        RECT 58.425 69.315 58.595 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_169/VNB
  PIN sky130_fd_sc_hd__decap_3_30/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 69.315 55.835 69.485 ;
    END
  END sky130_fd_sc_hd__decap_3_30/VNB
  PIN sky130_fd_sc_hd__buf_1_0/X
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 61.985 70.475 62.315 70.725 ;
        RECT 62.515 70.455 62.850 70.725 ;
        RECT 57.935 68.640 58.195 69.145 ;
        RECT 58.015 67.840 58.195 68.640 ;
        RECT 64.805 68.075 65.565 68.325 ;
        RECT 57.925 66.935 58.195 67.840 ;
      LAYER mcon ;
        RECT 62.105 70.505 62.275 70.675 ;
        RECT 62.565 70.505 62.735 70.675 ;
        RECT 57.965 68.805 58.135 68.975 ;
        RECT 64.865 68.125 65.035 68.295 ;
      LAYER met1 ;
        RECT 62.030 70.660 62.350 70.720 ;
        RECT 62.505 70.660 62.795 70.705 ;
        RECT 62.030 70.520 62.795 70.660 ;
        RECT 62.030 70.460 62.350 70.520 ;
        RECT 62.505 70.475 62.795 70.520 ;
        RECT 57.905 68.960 58.195 69.005 ;
        RECT 62.030 68.960 62.350 69.020 ;
        RECT 57.905 68.820 62.350 68.960 ;
        RECT 57.905 68.775 58.195 68.820 ;
        RECT 62.030 68.760 62.350 68.820 ;
        RECT 62.120 68.280 62.260 68.760 ;
        RECT 64.805 68.280 65.095 68.325 ;
        RECT 62.120 68.140 65.095 68.280 ;
        RECT 64.805 68.095 65.095 68.140 ;
      LAYER via ;
        RECT 62.060 70.460 62.320 70.720 ;
        RECT 62.060 68.760 62.320 69.020 ;
      LAYER met2 ;
        RECT 62.060 70.430 62.320 70.750 ;
        RECT 62.120 69.050 62.260 70.430 ;
        RECT 62.060 68.730 62.320 69.050 ;
    END
  END sky130_fd_sc_hd__buf_1_0/X
  PIN sky130_fd_sc_hd__buf_1_0/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 69.315 57.225 69.485 ;
    END
  END sky130_fd_sc_hd__buf_1_0/VNB
  PIN sky130_fd_sc_hd__fill_2_2/VNB
    PORT
      LAYER pwell ;
        RECT 63.955 69.340 64.115 69.450 ;
    END
  END sky130_fd_sc_hd__fill_2_2/VNB
  PIN sky130_fd_sc_hd__nand2_2_0/VNB
    PORT
      LAYER pwell ;
        RECT 64.870 69.315 65.040 69.485 ;
    END
  END sky130_fd_sc_hd__nand2_2_0/VNB
  PIN sky130_fd_sc_hd__ebufn_2_0/VNB
    PORT
      LAYER pwell ;
        RECT 67.160 69.315 67.340 69.485 ;
    END
  END sky130_fd_sc_hd__ebufn_2_0/VNB
  PIN sky130_ef_sc_hd__decap_12_168/VNB
    PORT
      LAYER pwell ;
        RECT 71.305 69.315 71.475 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_168/VNB
  PIN sky130_fd_sc_hd__decap_8_8/VNB
    PORT
      LAYER pwell ;
        RECT 76.825 69.315 76.995 69.485 ;
    END
  END sky130_fd_sc_hd__decap_8_8/VNB
  PIN sky130_fd_sc_hd__fill_2_1/VNB
    PORT
      LAYER pwell ;
        RECT 80.515 69.340 80.675 69.450 ;
    END
  END sky130_fd_sc_hd__fill_2_1/VNB
  PIN sky130_ef_sc_hd__decap_12_167/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 69.315 82.055 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_167/VNB
  PIN sky130_ef_sc_hd__decap_12_166/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 69.315 87.575 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_166/VNB
  PIN sky130_ef_sc_hd__decap_12_165/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 69.315 93.095 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_165/VNB
  PIN sky130_ef_sc_hd__decap_12_164/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 69.315 98.615 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_164/VNB
  PIN sky130_fd_sc_hd__decap_6_23/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 69.315 104.135 69.485 ;
    END
  END sky130_fd_sc_hd__decap_6_23/VNB
  PIN sky130_fd_sc_hd__fill_1_49/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 69.345 106.840 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_49/VNB
  PIN sky130_ef_sc_hd__decap_12_163/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 69.315 107.815 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_163/VNB
  PIN sky130_ef_sc_hd__decap_12_162/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 69.315 113.335 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_162/VNB
  PIN sky130_ef_sc_hd__decap_12_161/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 69.315 118.855 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_161/VNB
  PIN sky130_ef_sc_hd__decap_12_160/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 69.315 124.375 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_160/VNB
  PIN sky130_fd_sc_hd__decap_6_22/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 69.315 129.895 69.485 ;
    END
  END sky130_fd_sc_hd__decap_6_22/VNB
  PIN sky130_fd_sc_hd__fill_1_48/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 69.345 132.600 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_48/VNB
  PIN sky130_ef_sc_hd__decap_12_159/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 69.315 133.575 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_159/VNB
  PIN sky130_fd_sc_hd__decap_8_7/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 69.315 139.095 69.485 ;
    END
  END sky130_fd_sc_hd__decap_8_7/VNB
  PIN sky130_fd_sc_hd__fill_1_47/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 69.345 142.720 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_47/VNB
  PIN sky130_fd_sc_hd__decap_3_29/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 69.315 144.155 69.485 ;
    END
  END sky130_fd_sc_hd__decap_3_29/VNB
  PIN sky130_fd_sc_hd__fill_1_46/VNB
    PORT
      LAYER pwell ;
        RECT 60.720 69.345 60.840 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_46/VNB
  PIN sky130_fd_sc_hd__inv_2_1/Y
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 61.565 70.885 61.895 71.865 ;
        RECT 61.565 70.285 61.815 70.885 ;
        RECT 61.565 69.655 61.895 70.285 ;
    END
  END sky130_fd_sc_hd__inv_2_1/Y
  PIN sky130_fd_sc_hd__inv_2_1/VNB
    PORT
      LAYER pwell ;
        RECT 62.105 69.315 62.275 69.485 ;
    END
  END sky130_fd_sc_hd__inv_2_1/VNB
  PIN sky130_fd_sc_hd__nand2_1_0/Y
    ANTENNAGATEAREA 0.309000 ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 62.955 70.885 63.285 71.865 ;
        RECT 63.020 70.845 63.195 70.885 ;
        RECT 63.020 70.285 63.190 70.845 ;
        RECT 66.240 70.475 66.570 71.030 ;
        RECT 63.020 69.655 63.715 70.285 ;
      LAYER mcon ;
        RECT 63.025 70.845 63.195 71.015 ;
        RECT 66.245 70.845 66.415 71.015 ;
      LAYER met1 ;
        RECT 62.965 71.000 63.255 71.045 ;
        RECT 66.185 71.000 66.475 71.045 ;
        RECT 62.965 70.860 66.475 71.000 ;
        RECT 62.965 70.815 63.255 70.860 ;
        RECT 66.185 70.815 66.475 70.860 ;
    END
  END sky130_fd_sc_hd__nand2_1_0/Y
  PIN sky130_fd_sc_hd__nand2_1_0/VNB
    PORT
      LAYER pwell ;
        RECT 62.560 69.315 62.730 69.485 ;
    END
  END sky130_fd_sc_hd__nand2_1_0/VNB
  PIN sky130_fd_sc_hd__fill_2_0/VNB
    PORT
      LAYER pwell ;
        RECT 67.635 69.350 67.795 69.460 ;
    END
  END sky130_fd_sc_hd__fill_2_0/VNB
  PIN sky130_ef_sc_hd__decap_12_158/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 69.315 69.175 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_158/VNB
  PIN sky130_ef_sc_hd__decap_12_157/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 69.315 74.695 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_157/VNB
  PIN sky130_ef_sc_hd__decap_12_156/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 69.315 80.215 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_156/VNB
  PIN sky130_ef_sc_hd__decap_12_155/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 69.315 85.735 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_155/VNB
  PIN sky130_fd_sc_hd__decap_6_21/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 69.315 91.255 69.485 ;
    END
  END sky130_fd_sc_hd__decap_6_21/VNB
  PIN sky130_fd_sc_hd__fill_1_45/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 69.345 93.960 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_45/VNB
  PIN sky130_ef_sc_hd__decap_12_154/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 69.315 94.935 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_154/VNB
  PIN sky130_ef_sc_hd__decap_12_153/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 69.315 100.455 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_153/VNB
  PIN sky130_ef_sc_hd__decap_12_152/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 69.315 105.975 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_152/VNB
  PIN sky130_ef_sc_hd__decap_12_151/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 69.315 111.495 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_151/VNB
  PIN sky130_fd_sc_hd__decap_6_20/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 69.315 117.015 69.485 ;
    END
  END sky130_fd_sc_hd__decap_6_20/VNB
  PIN sky130_fd_sc_hd__fill_1_44/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 69.345 119.720 69.455 ;
    END
  END sky130_fd_sc_hd__fill_1_44/VNB
  PIN sky130_ef_sc_hd__decap_12_150/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 69.315 120.695 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_150/VNB
  PIN sky130_ef_sc_hd__decap_12_149/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 69.315 126.215 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_149/VNB
  PIN sky130_ef_sc_hd__decap_12_148/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 69.315 131.735 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_148/VNB
  PIN sky130_ef_sc_hd__decap_12_147/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 69.315 137.255 69.485 ;
    END
  END sky130_ef_sc_hd__decap_12_147/VNB
  PIN sky130_ef_sc_hd__decap_12_146/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 74.755 57.215 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_146/VNB
  PIN sky130_fd_sc_hd__decap_3_26/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 74.755 55.835 74.925 ;
    END
  END sky130_fd_sc_hd__decap_3_26/VNB
  PIN sky130_ef_sc_hd__decap_12_145/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 74.755 62.735 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_145/VNB
  PIN sky130_fd_sc_hd__decap_4_5/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 74.895 68.255 74.925 ;
        RECT 68.080 74.785 68.255 74.895 ;
        RECT 68.085 74.755 68.255 74.785 ;
    END
  END sky130_fd_sc_hd__decap_4_5/VNB
  PIN sky130_fd_sc_hd__fill_1_42/VNB
    PORT
      LAYER pwell ;
        RECT 69.920 74.785 70.040 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_42/VNB
  PIN sky130_fd_sc_hd__inv_2_0/Y
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 70.765 73.955 71.095 74.585 ;
        RECT 70.845 73.355 71.095 73.955 ;
        RECT 71.705 73.485 72.060 73.855 ;
        RECT 70.765 72.375 71.095 73.355 ;
      LAYER mcon ;
        RECT 70.845 73.565 71.015 73.735 ;
        RECT 71.765 73.565 71.935 73.735 ;
      LAYER met1 ;
        RECT 70.785 73.720 71.075 73.765 ;
        RECT 71.705 73.720 71.995 73.765 ;
        RECT 70.785 73.580 71.995 73.720 ;
        RECT 70.785 73.535 71.075 73.580 ;
        RECT 71.705 73.535 71.995 73.580 ;
    END
  END sky130_fd_sc_hd__inv_2_0/Y
  PIN sky130_fd_sc_hd__inv_2_0/VNB
    PORT
      LAYER pwell ;
        RECT 70.385 74.755 70.555 74.925 ;
    END
  END sky130_fd_sc_hd__inv_2_0/VNB
  PIN sky130_fd_sc_hd__buf_2_0/X
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 72.680 74.010 72.935 74.585 ;
        RECT 72.765 73.280 72.935 74.010 ;
        RECT 72.680 72.375 72.935 73.280 ;
    END
  END sky130_fd_sc_hd__buf_2_0/X
  PIN sky130_fd_sc_hd__buf_2_0/VNB
    PORT
      LAYER pwell ;
        RECT 71.765 74.755 71.935 74.925 ;
    END
  END sky130_fd_sc_hd__buf_2_0/VNB
  PIN sky130_ef_sc_hd__decap_12_144/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 74.755 73.775 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_144/VNB
  PIN sky130_fd_sc_hd__decap_4_4/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 74.755 79.295 74.925 ;
    END
  END sky130_fd_sc_hd__decap_4_4/VNB
  PIN sky130_fd_sc_hd__fill_1_41/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 74.785 81.080 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_41/VNB
  PIN sky130_ef_sc_hd__decap_12_143/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 74.755 82.055 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_143/VNB
  PIN sky130_ef_sc_hd__decap_12_142/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 74.755 87.575 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_142/VNB
  PIN sky130_ef_sc_hd__decap_12_141/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 74.755 93.095 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_141/VNB
  PIN sky130_ef_sc_hd__decap_12_140/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 74.755 98.615 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_140/VNB
  PIN sky130_fd_sc_hd__decap_6_19/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 74.755 104.135 74.925 ;
    END
  END sky130_fd_sc_hd__decap_6_19/VNB
  PIN sky130_fd_sc_hd__fill_1_40/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 74.785 106.840 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_40/VNB
  PIN sky130_ef_sc_hd__decap_12_139/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 74.755 107.815 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_139/VNB
  PIN sky130_ef_sc_hd__decap_12_138/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 74.755 113.335 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_138/VNB
  PIN sky130_ef_sc_hd__decap_12_137/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 74.755 118.855 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_137/VNB
  PIN sky130_ef_sc_hd__decap_12_136/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 74.755 124.375 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_136/VNB
  PIN sky130_fd_sc_hd__decap_6_18/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 74.755 129.895 74.925 ;
    END
  END sky130_fd_sc_hd__decap_6_18/VNB
  PIN sky130_fd_sc_hd__fill_1_39/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 74.785 132.600 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_39/VNB
  PIN sky130_ef_sc_hd__decap_12_135/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 74.755 133.575 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_135/VNB
  PIN sky130_fd_sc_hd__decap_8_5/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 74.755 139.095 74.925 ;
    END
  END sky130_fd_sc_hd__decap_8_5/VNB
  PIN sky130_fd_sc_hd__fill_1_38/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 74.785 142.720 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_38/VNB
  PIN sky130_fd_sc_hd__decap_3_25/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 74.755 144.155 74.925 ;
    END
  END sky130_fd_sc_hd__decap_3_25/VNB
  PIN sky130_ef_sc_hd__decap_12_132/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 74.755 69.175 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_132/VNB
  PIN sky130_ef_sc_hd__decap_12_131/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 74.755 74.695 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_131/VNB
  PIN sky130_ef_sc_hd__decap_12_130/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 74.755 80.215 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_130/VNB
  PIN sky130_ef_sc_hd__decap_12_129/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 74.755 85.735 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_129/VNB
  PIN sky130_fd_sc_hd__decap_6_17/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 74.755 91.255 74.925 ;
    END
  END sky130_fd_sc_hd__decap_6_17/VNB
  PIN sky130_fd_sc_hd__fill_1_36/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 74.785 93.960 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_36/VNB
  PIN sky130_ef_sc_hd__decap_12_128/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 74.755 94.935 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_128/VNB
  PIN sky130_ef_sc_hd__decap_12_127/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 74.755 100.455 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_127/VNB
  PIN sky130_ef_sc_hd__decap_12_126/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 74.755 105.975 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_126/VNB
  PIN sky130_ef_sc_hd__decap_12_125/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 74.755 111.495 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_125/VNB
  PIN sky130_fd_sc_hd__decap_6_16/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 74.755 117.015 74.925 ;
    END
  END sky130_fd_sc_hd__decap_6_16/VNB
  PIN sky130_fd_sc_hd__fill_1_35/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 74.785 119.720 74.895 ;
    END
  END sky130_fd_sc_hd__fill_1_35/VNB
  PIN sky130_ef_sc_hd__decap_12_124/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 74.755 120.695 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_124/VNB
  PIN sky130_ef_sc_hd__decap_12_123/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 74.755 126.215 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_123/VNB
  PIN sky130_ef_sc_hd__decap_12_122/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 74.755 131.735 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_122/VNB
  PIN sky130_ef_sc_hd__decap_12_121/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 74.755 137.255 74.925 ;
    END
  END sky130_ef_sc_hd__decap_12_121/VNB
  PIN sky130_ef_sc_hd__decap_12_120/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 80.195 57.215 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_120/VNB
  PIN sky130_fd_sc_hd__decap_3_22/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 80.195 55.835 80.365 ;
    END
  END sky130_fd_sc_hd__decap_3_22/VNB
  PIN sky130_ef_sc_hd__decap_12_118/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 80.195 62.735 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_118/VNB
  PIN sky130_ef_sc_hd__decap_12_116/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 80.335 68.255 80.365 ;
        RECT 68.080 80.225 68.255 80.335 ;
        RECT 68.085 80.195 68.255 80.225 ;
    END
  END sky130_ef_sc_hd__decap_12_116/VNB
  PIN sky130_ef_sc_hd__decap_12_115/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 80.195 69.175 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_115/VNB
  PIN sky130_ef_sc_hd__decap_12_114/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 80.195 73.775 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_114/VNB
  PIN sky130_fd_sc_hd__decap_4_3/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 80.195 79.295 80.365 ;
    END
  END sky130_fd_sc_hd__decap_4_3/VNB
  PIN sky130_ef_sc_hd__decap_12_113/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 80.195 74.695 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_113/VNB
  PIN sky130_fd_sc_hd__fill_1_32/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 80.225 81.080 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_32/VNB
  PIN sky130_ef_sc_hd__decap_12_112/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 80.195 82.055 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_112/VNB
  PIN sky130_ef_sc_hd__decap_12_111/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 80.195 80.215 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_111/VNB
  PIN sky130_ef_sc_hd__decap_12_110/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 80.195 87.575 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_110/VNB
  PIN sky130_ef_sc_hd__decap_12_109/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 80.195 85.735 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_109/VNB
  PIN sky130_fd_sc_hd__decap_6_15/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 80.195 91.255 80.365 ;
    END
  END sky130_fd_sc_hd__decap_6_15/VNB
  PIN sky130_ef_sc_hd__decap_12_108/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 80.195 93.095 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_108/VNB
  PIN sky130_fd_sc_hd__fill_1_31/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 80.225 93.960 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_31/VNB
  PIN sky130_ef_sc_hd__decap_12_107/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 80.195 94.935 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_107/VNB
  PIN sky130_ef_sc_hd__decap_12_106/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 80.195 98.615 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_106/VNB
  PIN sky130_ef_sc_hd__decap_12_105/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 80.195 100.455 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_105/VNB
  PIN sky130_fd_sc_hd__decap_6_14/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 80.195 104.135 80.365 ;
    END
  END sky130_fd_sc_hd__decap_6_14/VNB
  PIN sky130_fd_sc_hd__fill_1_30/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 80.225 106.840 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_30/VNB
  PIN sky130_ef_sc_hd__decap_12_104/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 80.195 107.815 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_104/VNB
  PIN sky130_ef_sc_hd__decap_12_103/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 80.195 105.975 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_103/VNB
  PIN sky130_ef_sc_hd__decap_12_102/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 80.195 113.335 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_102/VNB
  PIN sky130_ef_sc_hd__decap_12_101/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 80.195 111.495 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_101/VNB
  PIN sky130_ef_sc_hd__decap_12_100/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 80.195 118.855 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_100/VNB
  PIN sky130_fd_sc_hd__decap_6_13/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 80.195 117.015 80.365 ;
    END
  END sky130_fd_sc_hd__decap_6_13/VNB
  PIN sky130_fd_sc_hd__fill_1_29/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 80.225 119.720 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_29/VNB
  PIN sky130_ef_sc_hd__decap_12_99/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 80.195 120.695 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_99/VNB
  PIN sky130_ef_sc_hd__decap_12_98/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 80.195 124.375 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_98/VNB
  PIN sky130_ef_sc_hd__decap_12_97/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 80.195 126.215 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_97/VNB
  PIN sky130_fd_sc_hd__decap_6_12/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 80.195 129.895 80.365 ;
    END
  END sky130_fd_sc_hd__decap_6_12/VNB
  PIN sky130_ef_sc_hd__decap_12_96/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 80.195 131.735 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_96/VNB
  PIN sky130_fd_sc_hd__fill_1_28/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 80.225 132.600 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_28/VNB
  PIN sky130_ef_sc_hd__decap_12_95/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 80.195 133.575 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_95/VNB
  PIN sky130_ef_sc_hd__decap_12_94/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 80.195 137.255 80.365 ;
    END
  END sky130_ef_sc_hd__decap_12_94/VNB
  PIN sky130_fd_sc_hd__decap_8_4/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 80.195 139.095 80.365 ;
    END
  END sky130_fd_sc_hd__decap_8_4/VNB
  PIN sky130_fd_sc_hd__fill_1_27/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 80.225 142.720 80.335 ;
    END
  END sky130_fd_sc_hd__fill_1_27/VNB
  PIN sky130_fd_sc_hd__decap_3_20/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 80.195 144.155 80.365 ;
    END
  END sky130_fd_sc_hd__decap_3_20/VNB
  PIN sky130_ef_sc_hd__decap_12_93/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 85.635 57.215 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_93/VNB
  PIN sky130_fd_sc_hd__decap_3_18/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 85.635 55.835 85.805 ;
    END
  END sky130_fd_sc_hd__decap_3_18/VNB
  PIN sky130_ef_sc_hd__decap_12_92/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 85.635 62.735 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_92/VNB
  PIN sky130_ef_sc_hd__decap_12_91/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 85.775 68.255 85.805 ;
        RECT 68.080 85.665 68.255 85.775 ;
        RECT 68.085 85.635 68.255 85.665 ;
    END
  END sky130_ef_sc_hd__decap_12_91/VNB
  PIN sky130_ef_sc_hd__decap_12_90/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 85.635 73.775 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_90/VNB
  PIN sky130_fd_sc_hd__decap_4_2/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 85.635 79.295 85.805 ;
    END
  END sky130_fd_sc_hd__decap_4_2/VNB
  PIN sky130_fd_sc_hd__fill_1_25/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 85.665 81.080 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_25/VNB
  PIN sky130_ef_sc_hd__decap_12_89/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 85.635 82.055 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_89/VNB
  PIN sky130_ef_sc_hd__decap_12_88/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 85.635 87.575 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_88/VNB
  PIN sky130_ef_sc_hd__decap_12_87/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 85.635 93.095 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_87/VNB
  PIN sky130_ef_sc_hd__decap_12_86/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 85.635 98.615 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_86/VNB
  PIN sky130_fd_sc_hd__decap_6_11/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 85.635 104.135 85.805 ;
    END
  END sky130_fd_sc_hd__decap_6_11/VNB
  PIN sky130_fd_sc_hd__fill_1_24/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 85.665 106.840 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_24/VNB
  PIN sky130_ef_sc_hd__decap_12_85/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 85.635 107.815 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_85/VNB
  PIN sky130_ef_sc_hd__decap_12_84/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 85.635 113.335 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_84/VNB
  PIN sky130_ef_sc_hd__decap_12_83/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 85.635 118.855 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_83/VNB
  PIN sky130_ef_sc_hd__decap_12_82/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 85.635 124.375 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_82/VNB
  PIN sky130_fd_sc_hd__decap_6_10/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 85.635 129.895 85.805 ;
    END
  END sky130_fd_sc_hd__decap_6_10/VNB
  PIN sky130_fd_sc_hd__fill_1_23/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 85.665 132.600 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_23/VNB
  PIN sky130_ef_sc_hd__decap_12_81/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 85.635 133.575 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_81/VNB
  PIN sky130_fd_sc_hd__decap_8_3/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 85.635 139.095 85.805 ;
    END
  END sky130_fd_sc_hd__decap_8_3/VNB
  PIN sky130_fd_sc_hd__fill_1_22/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 85.665 142.720 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_22/VNB
  PIN sky130_fd_sc_hd__decap_3_17/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 85.635 144.155 85.805 ;
    END
  END sky130_fd_sc_hd__decap_3_17/VNB
  PIN sky130_ef_sc_hd__decap_12_78/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 85.635 69.175 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_78/VNB
  PIN sky130_ef_sc_hd__decap_12_77/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 85.635 74.695 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_77/VNB
  PIN sky130_ef_sc_hd__decap_12_76/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 85.635 80.215 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_76/VNB
  PIN sky130_ef_sc_hd__decap_12_75/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 85.635 85.735 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_75/VNB
  PIN sky130_fd_sc_hd__decap_6_9/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 85.635 91.255 85.805 ;
    END
  END sky130_fd_sc_hd__decap_6_9/VNB
  PIN sky130_fd_sc_hd__fill_1_20/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 85.665 93.960 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_20/VNB
  PIN sky130_ef_sc_hd__decap_12_74/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 85.635 94.935 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_74/VNB
  PIN sky130_ef_sc_hd__decap_12_73/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 85.635 100.455 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_73/VNB
  PIN sky130_ef_sc_hd__decap_12_72/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 85.635 105.975 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_72/VNB
  PIN sky130_ef_sc_hd__decap_12_71/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 85.635 111.495 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_71/VNB
  PIN sky130_fd_sc_hd__decap_6_8/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 85.635 117.015 85.805 ;
    END
  END sky130_fd_sc_hd__decap_6_8/VNB
  PIN sky130_fd_sc_hd__fill_1_19/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 85.665 119.720 85.775 ;
    END
  END sky130_fd_sc_hd__fill_1_19/VNB
  PIN sky130_ef_sc_hd__decap_12_70/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 85.635 120.695 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_70/VNB
  PIN sky130_ef_sc_hd__decap_12_69/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 85.635 126.215 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_69/VNB
  PIN sky130_ef_sc_hd__decap_12_68/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 85.635 131.735 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_68/VNB
  PIN sky130_ef_sc_hd__decap_12_67/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 85.635 137.255 85.805 ;
    END
  END sky130_ef_sc_hd__decap_12_67/VNB
  PIN sky130_ef_sc_hd__decap_12_66/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 91.075 57.215 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_66/VNB
  PIN sky130_fd_sc_hd__decap_3_14/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 91.075 55.835 91.245 ;
    END
  END sky130_fd_sc_hd__decap_3_14/VNB
  PIN sky130_ef_sc_hd__decap_12_65/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 91.075 62.735 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_65/VNB
  PIN sky130_ef_sc_hd__decap_12_64/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 91.215 68.255 91.245 ;
        RECT 68.080 91.105 68.255 91.215 ;
        RECT 68.085 91.075 68.255 91.105 ;
    END
  END sky130_ef_sc_hd__decap_12_64/VNB
  PIN sky130_ef_sc_hd__decap_12_63/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 91.075 73.775 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_63/VNB
  PIN sky130_fd_sc_hd__decap_4_1/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 91.075 79.295 91.245 ;
    END
  END sky130_fd_sc_hd__decap_4_1/VNB
  PIN sky130_fd_sc_hd__fill_1_17/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 91.105 81.080 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_17/VNB
  PIN sky130_ef_sc_hd__decap_12_62/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 91.075 82.055 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_62/VNB
  PIN sky130_ef_sc_hd__decap_12_61/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 91.075 87.575 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_61/VNB
  PIN sky130_ef_sc_hd__decap_12_60/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 91.075 93.095 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_60/VNB
  PIN sky130_ef_sc_hd__decap_12_59/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 91.075 98.615 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_59/VNB
  PIN sky130_fd_sc_hd__decap_6_7/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 91.075 104.135 91.245 ;
    END
  END sky130_fd_sc_hd__decap_6_7/VNB
  PIN sky130_fd_sc_hd__fill_1_16/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 91.105 106.840 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_16/VNB
  PIN sky130_ef_sc_hd__decap_12_58/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 91.075 107.815 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_58/VNB
  PIN sky130_ef_sc_hd__decap_12_57/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 91.075 113.335 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_57/VNB
  PIN sky130_ef_sc_hd__decap_12_56/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 91.075 118.855 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_56/VNB
  PIN sky130_ef_sc_hd__decap_12_55/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 91.075 124.375 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_55/VNB
  PIN sky130_fd_sc_hd__decap_6_6/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 91.075 129.895 91.245 ;
    END
  END sky130_fd_sc_hd__decap_6_6/VNB
  PIN sky130_fd_sc_hd__fill_1_15/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 91.105 132.600 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_15/VNB
  PIN sky130_ef_sc_hd__decap_12_54/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 91.075 133.575 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_54/VNB
  PIN sky130_fd_sc_hd__decap_8_2/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 91.075 139.095 91.245 ;
    END
  END sky130_fd_sc_hd__decap_8_2/VNB
  PIN sky130_fd_sc_hd__fill_1_14/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 91.105 142.720 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_14/VNB
  PIN sky130_fd_sc_hd__decap_3_13/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 91.075 144.155 91.245 ;
    END
  END sky130_fd_sc_hd__decap_3_13/VNB
  PIN sky130_ef_sc_hd__decap_12_51/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 91.075 69.175 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_51/VNB
  PIN sky130_ef_sc_hd__decap_12_50/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 91.075 74.695 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_50/VNB
  PIN sky130_ef_sc_hd__decap_12_49/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 91.075 80.215 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_49/VNB
  PIN sky130_ef_sc_hd__decap_12_48/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 91.075 85.735 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_48/VNB
  PIN sky130_fd_sc_hd__decap_6_5/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 91.075 91.255 91.245 ;
    END
  END sky130_fd_sc_hd__decap_6_5/VNB
  PIN sky130_fd_sc_hd__fill_1_12/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 91.105 93.960 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_12/VNB
  PIN sky130_ef_sc_hd__decap_12_47/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 91.075 94.935 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_47/VNB
  PIN sky130_ef_sc_hd__decap_12_46/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 91.075 100.455 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_46/VNB
  PIN sky130_ef_sc_hd__decap_12_45/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 91.075 105.975 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_45/VNB
  PIN sky130_ef_sc_hd__decap_12_44/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 91.075 111.495 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_44/VNB
  PIN sky130_fd_sc_hd__decap_6_4/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 91.075 117.015 91.245 ;
    END
  END sky130_fd_sc_hd__decap_6_4/VNB
  PIN sky130_fd_sc_hd__fill_1_11/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 91.105 119.720 91.215 ;
    END
  END sky130_fd_sc_hd__fill_1_11/VNB
  PIN sky130_ef_sc_hd__decap_12_43/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 91.075 120.695 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_43/VNB
  PIN sky130_ef_sc_hd__decap_12_42/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 91.075 126.215 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_42/VNB
  PIN sky130_ef_sc_hd__decap_12_41/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 91.075 131.735 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_41/VNB
  PIN sky130_ef_sc_hd__decap_12_40/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 91.075 137.255 91.245 ;
    END
  END sky130_ef_sc_hd__decap_12_40/VNB
  PIN sky130_ef_sc_hd__decap_12_39/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 96.515 57.215 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_39/VNB
  PIN sky130_fd_sc_hd__decap_3_10/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 96.515 55.835 96.685 ;
    END
  END sky130_fd_sc_hd__decap_3_10/VNB
  PIN sky130_ef_sc_hd__decap_12_38/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 96.515 62.735 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_38/VNB
  PIN sky130_ef_sc_hd__decap_12_37/VNB
    PORT
      LAYER pwell ;
        RECT 68.085 96.655 68.255 96.685 ;
        RECT 68.080 96.545 68.255 96.655 ;
        RECT 68.085 96.515 68.255 96.545 ;
    END
  END sky130_ef_sc_hd__decap_12_37/VNB
  PIN sky130_ef_sc_hd__decap_12_36/VNB
    PORT
      LAYER pwell ;
        RECT 73.605 96.515 73.775 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_36/VNB
  PIN sky130_fd_sc_hd__decap_4_0/VNB
    PORT
      LAYER pwell ;
        RECT 79.125 96.515 79.295 96.685 ;
    END
  END sky130_fd_sc_hd__decap_4_0/VNB
  PIN sky130_fd_sc_hd__fill_1_9/VNB
    PORT
      LAYER pwell ;
        RECT 80.960 96.545 81.080 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_9/VNB
  PIN sky130_ef_sc_hd__decap_12_35/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 96.515 82.055 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_35/VNB
  PIN sky130_ef_sc_hd__decap_12_34/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 96.515 87.575 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_34/VNB
  PIN sky130_ef_sc_hd__decap_12_33/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 96.515 93.095 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_33/VNB
  PIN sky130_ef_sc_hd__decap_12_32/VNB
    PORT
      LAYER pwell ;
        RECT 98.445 96.515 98.615 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_32/VNB
  PIN sky130_fd_sc_hd__decap_6_3/VNB
    PORT
      LAYER pwell ;
        RECT 103.965 96.515 104.135 96.685 ;
    END
  END sky130_fd_sc_hd__decap_6_3/VNB
  PIN sky130_fd_sc_hd__fill_1_8/VNB
    PORT
      LAYER pwell ;
        RECT 106.720 96.545 106.840 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_8/VNB
  PIN sky130_ef_sc_hd__decap_12_31/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 96.515 107.815 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_31/VNB
  PIN sky130_ef_sc_hd__decap_12_30/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 96.515 113.335 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_30/VNB
  PIN sky130_ef_sc_hd__decap_12_29/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 96.515 118.855 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_29/VNB
  PIN sky130_ef_sc_hd__decap_12_28/VNB
    PORT
      LAYER pwell ;
        RECT 124.205 96.515 124.375 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_28/VNB
  PIN sky130_fd_sc_hd__decap_6_2/VNB
    PORT
      LAYER pwell ;
        RECT 129.725 96.515 129.895 96.685 ;
    END
  END sky130_fd_sc_hd__decap_6_2/VNB
  PIN sky130_fd_sc_hd__fill_1_7/VNB
    PORT
      LAYER pwell ;
        RECT 132.480 96.545 132.600 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_7/VNB
  PIN sky130_ef_sc_hd__decap_12_27/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 96.515 133.575 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_27/VNB
  PIN sky130_fd_sc_hd__decap_8_1/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 96.515 139.095 96.685 ;
    END
  END sky130_fd_sc_hd__decap_8_1/VNB
  PIN sky130_fd_sc_hd__fill_1_6/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 96.545 142.720 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_6/VNB
  PIN sky130_fd_sc_hd__decap_3_9/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 96.515 144.155 96.685 ;
    END
  END sky130_fd_sc_hd__decap_3_9/VNB
  PIN sky130_ef_sc_hd__decap_12_25/VNB
    PORT
      LAYER pwell ;
        RECT 57.045 101.955 57.215 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_25/VNB
  PIN sky130_fd_sc_hd__decap_3_7/VNB
    PORT
      LAYER pwell ;
        RECT 55.665 101.955 55.835 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_7/VNB
  PIN sky130_ef_sc_hd__decap_12_23/VNB
    PORT
      LAYER pwell ;
        RECT 62.565 101.955 62.735 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_23/VNB
  PIN sky130_ef_sc_hd__decap_12_22/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 96.515 69.175 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_22/VNB
  PIN sky130_fd_sc_hd__fill_1_4/VNB
    PORT
      LAYER pwell ;
        RECT 68.080 101.985 68.200 102.095 ;
    END
  END sky130_fd_sc_hd__fill_1_4/VNB
  PIN sky130_ef_sc_hd__decap_12_21/VNB
    PORT
      LAYER pwell ;
        RECT 69.005 101.955 69.175 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_21/VNB
  PIN sky130_ef_sc_hd__decap_12_20/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 96.515 74.695 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_20/VNB
  PIN sky130_ef_sc_hd__decap_12_19/VNB
    PORT
      LAYER pwell ;
        RECT 74.525 101.955 74.695 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_19/VNB
  PIN sky130_ef_sc_hd__decap_12_18/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 96.515 80.215 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_18/VNB
  PIN sky130_fd_sc_hd__decap_3_6/VNB
    PORT
      LAYER pwell ;
        RECT 80.045 101.955 80.215 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_6/VNB
  PIN sky130_ef_sc_hd__decap_12_17/VNB
    PORT
      LAYER pwell ;
        RECT 81.885 101.955 82.055 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_17/VNB
  PIN sky130_ef_sc_hd__decap_12_16/VNB
    PORT
      LAYER pwell ;
        RECT 85.565 96.515 85.735 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_16/VNB
  PIN sky130_fd_sc_hd__decap_6_1/VNB
    PORT
      LAYER pwell ;
        RECT 91.085 96.515 91.255 96.685 ;
    END
  END sky130_fd_sc_hd__decap_6_1/VNB
  PIN sky130_ef_sc_hd__decap_12_15/VNB
    PORT
      LAYER pwell ;
        RECT 87.405 101.955 87.575 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_15/VNB
  PIN sky130_fd_sc_hd__fill_1_3/VNB
    PORT
      LAYER pwell ;
        RECT 93.840 96.545 93.960 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_3/VNB
  PIN sky130_ef_sc_hd__decap_12_14/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 96.515 94.935 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_14/VNB
  PIN sky130_fd_sc_hd__decap_3_5/VNB
    PORT
      LAYER pwell ;
        RECT 92.925 101.955 93.095 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_5/VNB
  PIN sky130_ef_sc_hd__decap_12_13/VNB
    PORT
      LAYER pwell ;
        RECT 94.765 101.955 94.935 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_13/VNB
  PIN sky130_ef_sc_hd__decap_12_12/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 96.515 100.455 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_12/VNB
  PIN sky130_ef_sc_hd__decap_12_11/VNB
    PORT
      LAYER pwell ;
        RECT 100.285 101.955 100.455 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_11/VNB
  PIN sky130_ef_sc_hd__decap_12_10/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 96.515 105.975 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_10/VNB
  PIN sky130_fd_sc_hd__decap_3_4/VNB
    PORT
      LAYER pwell ;
        RECT 105.805 101.955 105.975 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_4/VNB
  PIN sky130_ef_sc_hd__decap_12_9/VNB
    PORT
      LAYER pwell ;
        RECT 107.645 101.955 107.815 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_9/VNB
  PIN sky130_ef_sc_hd__decap_12_8/VNB
    PORT
      LAYER pwell ;
        RECT 111.325 96.515 111.495 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_8/VNB
  PIN sky130_ef_sc_hd__decap_12_7/VNB
    PORT
      LAYER pwell ;
        RECT 113.165 101.955 113.335 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_7/VNB
  PIN sky130_fd_sc_hd__decap_6_0/VNB
    PORT
      LAYER pwell ;
        RECT 116.845 96.515 117.015 96.685 ;
    END
  END sky130_fd_sc_hd__decap_6_0/VNB
  PIN sky130_fd_sc_hd__fill_1_2/VNB
    PORT
      LAYER pwell ;
        RECT 119.600 96.545 119.720 96.655 ;
    END
  END sky130_fd_sc_hd__fill_1_2/VNB
  PIN sky130_ef_sc_hd__decap_12_6/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 96.515 120.695 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_6/VNB
  PIN sky130_fd_sc_hd__decap_3_3/VNB
    PORT
      LAYER pwell ;
        RECT 118.685 101.955 118.855 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_3/VNB
  PIN sky130_ef_sc_hd__decap_12_5/VNB
    PORT
      LAYER pwell ;
        RECT 120.525 101.955 120.695 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_5/VNB
  PIN sky130_ef_sc_hd__decap_12_4/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 96.515 126.215 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_4/VNB
  PIN sky130_ef_sc_hd__decap_12_3/VNB
    PORT
      LAYER pwell ;
        RECT 126.045 101.955 126.215 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_3/VNB
  PIN sky130_ef_sc_hd__decap_12_2/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 96.515 131.735 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_2/VNB
  PIN sky130_fd_sc_hd__decap_3_2/VNB
    PORT
      LAYER pwell ;
        RECT 131.565 101.955 131.735 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_2/VNB
  PIN sky130_ef_sc_hd__decap_12_1/VNB
    PORT
      LAYER pwell ;
        RECT 137.085 96.515 137.255 96.685 ;
    END
  END sky130_ef_sc_hd__decap_12_1/VNB
  PIN sky130_ef_sc_hd__decap_12_0/VNB
    PORT
      LAYER pwell ;
        RECT 133.405 101.955 133.575 102.125 ;
    END
  END sky130_ef_sc_hd__decap_12_0/VNB
  PIN sky130_fd_sc_hd__decap_8_0/VNB
    PORT
      LAYER pwell ;
        RECT 138.925 101.955 139.095 102.125 ;
    END
  END sky130_fd_sc_hd__decap_8_0/VNB
  PIN sky130_fd_sc_hd__fill_1_0/VNB
    PORT
      LAYER pwell ;
        RECT 142.600 101.985 142.720 102.095 ;
    END
  END sky130_fd_sc_hd__fill_1_0/VNB
  PIN sky130_fd_sc_hd__decap_3_0/VNB
    PORT
      LAYER pwell ;
        RECT 143.985 101.955 144.155 102.125 ;
    END
  END sky130_fd_sc_hd__decap_3_0/VNB
  OBS
      LAYER li1 ;
        RECT 71.795 74.205 71.965 74.585 ;
        RECT 71.795 74.035 72.510 74.205 ;
        RECT 72.340 73.845 72.510 74.035 ;
        RECT 72.340 73.515 72.595 73.845 ;
        RECT 72.340 73.305 72.510 73.515 ;
        RECT 71.795 73.135 72.510 73.305 ;
        RECT 71.795 72.375 71.965 73.135 ;
        RECT 66.210 71.405 66.465 71.860 ;
        RECT 67.135 71.405 67.395 71.865 ;
        RECT 65.675 71.200 66.465 71.405 ;
        RECT 65.675 70.725 66.070 71.200 ;
        RECT 64.395 70.395 64.775 70.725 ;
        RECT 64.945 70.475 66.070 70.725 ;
        RECT 64.525 70.305 64.775 70.395 ;
        RECT 64.525 70.135 65.625 70.305 ;
        RECT 65.455 69.865 65.625 70.135 ;
        RECT 65.795 70.285 66.070 70.475 ;
        RECT 66.740 71.185 67.395 71.405 ;
        RECT 65.795 70.035 66.125 70.285 ;
        RECT 66.740 70.225 66.955 71.185 ;
        RECT 66.295 70.015 67.395 70.225 ;
        RECT 66.295 69.865 66.465 70.015 ;
        RECT 65.455 69.655 66.465 69.865 ;
        RECT 67.135 69.680 67.395 70.015 ;
        RECT 57.075 68.765 57.245 69.145 ;
        RECT 57.075 68.595 57.740 68.765 ;
        RECT 57.570 68.340 57.740 68.595 ;
        RECT 64.805 68.685 65.145 69.145 ;
        RECT 65.655 68.935 66.825 69.145 ;
        RECT 65.655 68.685 65.905 68.935 ;
        RECT 66.495 68.915 66.825 68.935 ;
        RECT 64.805 68.515 65.905 68.685 ;
        RECT 67.105 68.785 67.365 69.120 ;
        RECT 68.040 68.805 68.750 69.145 ;
        RECT 57.570 68.010 57.845 68.340 ;
        RECT 57.570 67.865 57.740 68.010 ;
        RECT 57.065 67.695 57.740 67.865 ;
        RECT 57.065 66.935 57.245 67.695 ;
        RECT 67.105 67.555 67.340 68.785 ;
        RECT 68.470 68.375 68.750 68.805 ;
        RECT 68.920 68.745 69.190 69.145 ;
        RECT 69.860 68.935 71.070 69.125 ;
        RECT 69.860 68.745 70.145 68.935 ;
        RECT 68.920 68.545 70.145 68.745 ;
        RECT 68.470 68.125 69.985 68.375 ;
        RECT 70.265 68.125 70.675 68.375 ;
        RECT 68.470 67.955 68.755 68.125 ;
        RECT 68.140 67.635 68.755 67.955 ;
        RECT 67.105 66.935 67.365 67.555 ;
        RECT 68.140 66.935 68.430 67.635 ;
        RECT 68.620 67.295 70.145 67.465 ;
        RECT 68.620 66.935 68.830 67.295 ;
        RECT 69.500 67.105 70.145 67.295 ;
        RECT 70.815 67.105 71.075 67.605 ;
        RECT 69.500 66.935 71.075 67.105 ;
        RECT 57.065 65.665 57.245 66.425 ;
        RECT 57.065 65.495 57.740 65.665 ;
        RECT 57.570 65.350 57.740 65.495 ;
        RECT 57.570 65.020 57.845 65.350 ;
        RECT 57.570 64.765 57.740 65.020 ;
        RECT 57.075 64.595 57.740 64.765 ;
        RECT 57.075 64.215 57.245 64.595 ;
        RECT 65.815 63.325 65.985 63.705 ;
        RECT 65.815 63.155 66.480 63.325 ;
        RECT 66.310 62.900 66.480 63.155 ;
        RECT 66.310 62.570 66.595 62.900 ;
        RECT 66.310 62.425 66.480 62.570 ;
        RECT 65.815 62.255 66.480 62.425 ;
        RECT 65.815 61.495 65.985 62.255 ;
        RECT 61.860 57.625 62.105 58.230 ;
        RECT 63.840 57.900 64.370 58.265 ;
        RECT 64.195 57.865 64.370 57.900 ;
        RECT 66.910 57.900 67.440 58.265 ;
        RECT 66.910 57.865 67.085 57.900 ;
        RECT 64.195 57.695 65.125 57.865 ;
        RECT 61.585 57.455 62.815 57.625 ;
        RECT 61.585 56.645 61.925 57.455 ;
        RECT 61.585 56.235 62.100 56.645 ;
        RECT 64.195 56.565 64.365 57.695 ;
        RECT 64.955 57.525 65.125 57.695 ;
        RECT 66.155 57.695 67.085 57.865 ;
        RECT 66.155 57.525 66.325 57.695 ;
        RECT 64.955 57.195 65.210 57.525 ;
        RECT 66.070 57.195 66.325 57.525 ;
        RECT 63.240 56.395 64.365 56.565 ;
        RECT 66.915 56.565 67.085 57.695 ;
        RECT 69.175 57.625 69.420 58.230 ;
        RECT 68.465 57.455 69.695 57.625 ;
        RECT 69.355 56.645 69.695 57.455 ;
        RECT 66.915 56.395 68.040 56.565 ;
        RECT 69.180 56.235 69.695 56.645 ;
        RECT 65.345 54.785 65.525 55.545 ;
        RECT 65.345 54.615 66.020 54.785 ;
        RECT 65.850 54.470 66.020 54.615 ;
        RECT 65.850 54.140 66.125 54.470 ;
        RECT 65.850 53.885 66.020 54.140 ;
        RECT 65.355 53.715 66.020 53.885 ;
        RECT 65.355 53.335 65.525 53.715 ;
      LAYER mcon ;
        RECT 67.170 68.125 67.340 68.295 ;
        RECT 70.400 68.125 70.570 68.295 ;
      LAYER met1 ;
        RECT 67.105 68.280 67.400 68.325 ;
        RECT 70.340 68.280 70.630 68.325 ;
        RECT 67.105 68.140 70.630 68.280 ;
        RECT 67.105 68.095 67.400 68.140 ;
        RECT 70.340 68.095 70.630 68.140 ;
  END
END dgiota
END LIBRARY

